magic
tech sky130A
magscale 1 2
timestamp 1697533315
<< nwell >>
rect -1809 -1597 1809 1597
<< mvpmos >>
rect -1551 -1300 -1451 1300
rect -1393 -1300 -1293 1300
rect -1235 -1300 -1135 1300
rect -1077 -1300 -977 1300
rect -919 -1300 -819 1300
rect -761 -1300 -661 1300
rect -603 -1300 -503 1300
rect -445 -1300 -345 1300
rect -287 -1300 -187 1300
rect -129 -1300 -29 1300
rect 29 -1300 129 1300
rect 187 -1300 287 1300
rect 345 -1300 445 1300
rect 503 -1300 603 1300
rect 661 -1300 761 1300
rect 819 -1300 919 1300
rect 977 -1300 1077 1300
rect 1135 -1300 1235 1300
rect 1293 -1300 1393 1300
rect 1451 -1300 1551 1300
<< mvpdiff >>
rect -1609 1288 -1551 1300
rect -1609 -1288 -1597 1288
rect -1563 -1288 -1551 1288
rect -1609 -1300 -1551 -1288
rect -1451 1288 -1393 1300
rect -1451 -1288 -1439 1288
rect -1405 -1288 -1393 1288
rect -1451 -1300 -1393 -1288
rect -1293 1288 -1235 1300
rect -1293 -1288 -1281 1288
rect -1247 -1288 -1235 1288
rect -1293 -1300 -1235 -1288
rect -1135 1288 -1077 1300
rect -1135 -1288 -1123 1288
rect -1089 -1288 -1077 1288
rect -1135 -1300 -1077 -1288
rect -977 1288 -919 1300
rect -977 -1288 -965 1288
rect -931 -1288 -919 1288
rect -977 -1300 -919 -1288
rect -819 1288 -761 1300
rect -819 -1288 -807 1288
rect -773 -1288 -761 1288
rect -819 -1300 -761 -1288
rect -661 1288 -603 1300
rect -661 -1288 -649 1288
rect -615 -1288 -603 1288
rect -661 -1300 -603 -1288
rect -503 1288 -445 1300
rect -503 -1288 -491 1288
rect -457 -1288 -445 1288
rect -503 -1300 -445 -1288
rect -345 1288 -287 1300
rect -345 -1288 -333 1288
rect -299 -1288 -287 1288
rect -345 -1300 -287 -1288
rect -187 1288 -129 1300
rect -187 -1288 -175 1288
rect -141 -1288 -129 1288
rect -187 -1300 -129 -1288
rect -29 1288 29 1300
rect -29 -1288 -17 1288
rect 17 -1288 29 1288
rect -29 -1300 29 -1288
rect 129 1288 187 1300
rect 129 -1288 141 1288
rect 175 -1288 187 1288
rect 129 -1300 187 -1288
rect 287 1288 345 1300
rect 287 -1288 299 1288
rect 333 -1288 345 1288
rect 287 -1300 345 -1288
rect 445 1288 503 1300
rect 445 -1288 457 1288
rect 491 -1288 503 1288
rect 445 -1300 503 -1288
rect 603 1288 661 1300
rect 603 -1288 615 1288
rect 649 -1288 661 1288
rect 603 -1300 661 -1288
rect 761 1288 819 1300
rect 761 -1288 773 1288
rect 807 -1288 819 1288
rect 761 -1300 819 -1288
rect 919 1288 977 1300
rect 919 -1288 931 1288
rect 965 -1288 977 1288
rect 919 -1300 977 -1288
rect 1077 1288 1135 1300
rect 1077 -1288 1089 1288
rect 1123 -1288 1135 1288
rect 1077 -1300 1135 -1288
rect 1235 1288 1293 1300
rect 1235 -1288 1247 1288
rect 1281 -1288 1293 1288
rect 1235 -1300 1293 -1288
rect 1393 1288 1451 1300
rect 1393 -1288 1405 1288
rect 1439 -1288 1451 1288
rect 1393 -1300 1451 -1288
rect 1551 1288 1609 1300
rect 1551 -1288 1563 1288
rect 1597 -1288 1609 1288
rect 1551 -1300 1609 -1288
<< mvpdiffc >>
rect -1597 -1288 -1563 1288
rect -1439 -1288 -1405 1288
rect -1281 -1288 -1247 1288
rect -1123 -1288 -1089 1288
rect -965 -1288 -931 1288
rect -807 -1288 -773 1288
rect -649 -1288 -615 1288
rect -491 -1288 -457 1288
rect -333 -1288 -299 1288
rect -175 -1288 -141 1288
rect -17 -1288 17 1288
rect 141 -1288 175 1288
rect 299 -1288 333 1288
rect 457 -1288 491 1288
rect 615 -1288 649 1288
rect 773 -1288 807 1288
rect 931 -1288 965 1288
rect 1089 -1288 1123 1288
rect 1247 -1288 1281 1288
rect 1405 -1288 1439 1288
rect 1563 -1288 1597 1288
<< mvnsubdiff >>
rect -1743 1519 1743 1531
rect -1743 1485 -1635 1519
rect 1635 1485 1743 1519
rect -1743 1473 1743 1485
rect -1743 1423 -1685 1473
rect -1743 -1423 -1731 1423
rect -1697 -1423 -1685 1423
rect 1685 1423 1743 1473
rect -1743 -1473 -1685 -1423
rect 1685 -1423 1697 1423
rect 1731 -1423 1743 1423
rect 1685 -1473 1743 -1423
rect -1743 -1485 1743 -1473
rect -1743 -1519 -1635 -1485
rect 1635 -1519 1743 -1485
rect -1743 -1531 1743 -1519
<< mvnsubdiffcont >>
rect -1635 1485 1635 1519
rect -1731 -1423 -1697 1423
rect 1697 -1423 1731 1423
rect -1635 -1519 1635 -1485
<< poly >>
rect -1551 1381 -1451 1397
rect -1551 1347 -1535 1381
rect -1467 1347 -1451 1381
rect -1551 1300 -1451 1347
rect -1393 1381 -1293 1397
rect -1393 1347 -1377 1381
rect -1309 1347 -1293 1381
rect -1393 1300 -1293 1347
rect -1235 1381 -1135 1397
rect -1235 1347 -1219 1381
rect -1151 1347 -1135 1381
rect -1235 1300 -1135 1347
rect -1077 1381 -977 1397
rect -1077 1347 -1061 1381
rect -993 1347 -977 1381
rect -1077 1300 -977 1347
rect -919 1381 -819 1397
rect -919 1347 -903 1381
rect -835 1347 -819 1381
rect -919 1300 -819 1347
rect -761 1381 -661 1397
rect -761 1347 -745 1381
rect -677 1347 -661 1381
rect -761 1300 -661 1347
rect -603 1381 -503 1397
rect -603 1347 -587 1381
rect -519 1347 -503 1381
rect -603 1300 -503 1347
rect -445 1381 -345 1397
rect -445 1347 -429 1381
rect -361 1347 -345 1381
rect -445 1300 -345 1347
rect -287 1381 -187 1397
rect -287 1347 -271 1381
rect -203 1347 -187 1381
rect -287 1300 -187 1347
rect -129 1381 -29 1397
rect -129 1347 -113 1381
rect -45 1347 -29 1381
rect -129 1300 -29 1347
rect 29 1381 129 1397
rect 29 1347 45 1381
rect 113 1347 129 1381
rect 29 1300 129 1347
rect 187 1381 287 1397
rect 187 1347 203 1381
rect 271 1347 287 1381
rect 187 1300 287 1347
rect 345 1381 445 1397
rect 345 1347 361 1381
rect 429 1347 445 1381
rect 345 1300 445 1347
rect 503 1381 603 1397
rect 503 1347 519 1381
rect 587 1347 603 1381
rect 503 1300 603 1347
rect 661 1381 761 1397
rect 661 1347 677 1381
rect 745 1347 761 1381
rect 661 1300 761 1347
rect 819 1381 919 1397
rect 819 1347 835 1381
rect 903 1347 919 1381
rect 819 1300 919 1347
rect 977 1381 1077 1397
rect 977 1347 993 1381
rect 1061 1347 1077 1381
rect 977 1300 1077 1347
rect 1135 1381 1235 1397
rect 1135 1347 1151 1381
rect 1219 1347 1235 1381
rect 1135 1300 1235 1347
rect 1293 1381 1393 1397
rect 1293 1347 1309 1381
rect 1377 1347 1393 1381
rect 1293 1300 1393 1347
rect 1451 1381 1551 1397
rect 1451 1347 1467 1381
rect 1535 1347 1551 1381
rect 1451 1300 1551 1347
rect -1551 -1347 -1451 -1300
rect -1551 -1381 -1535 -1347
rect -1467 -1381 -1451 -1347
rect -1551 -1397 -1451 -1381
rect -1393 -1347 -1293 -1300
rect -1393 -1381 -1377 -1347
rect -1309 -1381 -1293 -1347
rect -1393 -1397 -1293 -1381
rect -1235 -1347 -1135 -1300
rect -1235 -1381 -1219 -1347
rect -1151 -1381 -1135 -1347
rect -1235 -1397 -1135 -1381
rect -1077 -1347 -977 -1300
rect -1077 -1381 -1061 -1347
rect -993 -1381 -977 -1347
rect -1077 -1397 -977 -1381
rect -919 -1347 -819 -1300
rect -919 -1381 -903 -1347
rect -835 -1381 -819 -1347
rect -919 -1397 -819 -1381
rect -761 -1347 -661 -1300
rect -761 -1381 -745 -1347
rect -677 -1381 -661 -1347
rect -761 -1397 -661 -1381
rect -603 -1347 -503 -1300
rect -603 -1381 -587 -1347
rect -519 -1381 -503 -1347
rect -603 -1397 -503 -1381
rect -445 -1347 -345 -1300
rect -445 -1381 -429 -1347
rect -361 -1381 -345 -1347
rect -445 -1397 -345 -1381
rect -287 -1347 -187 -1300
rect -287 -1381 -271 -1347
rect -203 -1381 -187 -1347
rect -287 -1397 -187 -1381
rect -129 -1347 -29 -1300
rect -129 -1381 -113 -1347
rect -45 -1381 -29 -1347
rect -129 -1397 -29 -1381
rect 29 -1347 129 -1300
rect 29 -1381 45 -1347
rect 113 -1381 129 -1347
rect 29 -1397 129 -1381
rect 187 -1347 287 -1300
rect 187 -1381 203 -1347
rect 271 -1381 287 -1347
rect 187 -1397 287 -1381
rect 345 -1347 445 -1300
rect 345 -1381 361 -1347
rect 429 -1381 445 -1347
rect 345 -1397 445 -1381
rect 503 -1347 603 -1300
rect 503 -1381 519 -1347
rect 587 -1381 603 -1347
rect 503 -1397 603 -1381
rect 661 -1347 761 -1300
rect 661 -1381 677 -1347
rect 745 -1381 761 -1347
rect 661 -1397 761 -1381
rect 819 -1347 919 -1300
rect 819 -1381 835 -1347
rect 903 -1381 919 -1347
rect 819 -1397 919 -1381
rect 977 -1347 1077 -1300
rect 977 -1381 993 -1347
rect 1061 -1381 1077 -1347
rect 977 -1397 1077 -1381
rect 1135 -1347 1235 -1300
rect 1135 -1381 1151 -1347
rect 1219 -1381 1235 -1347
rect 1135 -1397 1235 -1381
rect 1293 -1347 1393 -1300
rect 1293 -1381 1309 -1347
rect 1377 -1381 1393 -1347
rect 1293 -1397 1393 -1381
rect 1451 -1347 1551 -1300
rect 1451 -1381 1467 -1347
rect 1535 -1381 1551 -1347
rect 1451 -1397 1551 -1381
<< polycont >>
rect -1535 1347 -1467 1381
rect -1377 1347 -1309 1381
rect -1219 1347 -1151 1381
rect -1061 1347 -993 1381
rect -903 1347 -835 1381
rect -745 1347 -677 1381
rect -587 1347 -519 1381
rect -429 1347 -361 1381
rect -271 1347 -203 1381
rect -113 1347 -45 1381
rect 45 1347 113 1381
rect 203 1347 271 1381
rect 361 1347 429 1381
rect 519 1347 587 1381
rect 677 1347 745 1381
rect 835 1347 903 1381
rect 993 1347 1061 1381
rect 1151 1347 1219 1381
rect 1309 1347 1377 1381
rect 1467 1347 1535 1381
rect -1535 -1381 -1467 -1347
rect -1377 -1381 -1309 -1347
rect -1219 -1381 -1151 -1347
rect -1061 -1381 -993 -1347
rect -903 -1381 -835 -1347
rect -745 -1381 -677 -1347
rect -587 -1381 -519 -1347
rect -429 -1381 -361 -1347
rect -271 -1381 -203 -1347
rect -113 -1381 -45 -1347
rect 45 -1381 113 -1347
rect 203 -1381 271 -1347
rect 361 -1381 429 -1347
rect 519 -1381 587 -1347
rect 677 -1381 745 -1347
rect 835 -1381 903 -1347
rect 993 -1381 1061 -1347
rect 1151 -1381 1219 -1347
rect 1309 -1381 1377 -1347
rect 1467 -1381 1535 -1347
<< locali >>
rect -1731 1485 -1635 1519
rect 1635 1485 1731 1519
rect -1731 1423 -1697 1485
rect 1697 1423 1731 1485
rect -1551 1347 -1535 1381
rect -1467 1347 -1451 1381
rect -1393 1347 -1377 1381
rect -1309 1347 -1293 1381
rect -1235 1347 -1219 1381
rect -1151 1347 -1135 1381
rect -1077 1347 -1061 1381
rect -993 1347 -977 1381
rect -919 1347 -903 1381
rect -835 1347 -819 1381
rect -761 1347 -745 1381
rect -677 1347 -661 1381
rect -603 1347 -587 1381
rect -519 1347 -503 1381
rect -445 1347 -429 1381
rect -361 1347 -345 1381
rect -287 1347 -271 1381
rect -203 1347 -187 1381
rect -129 1347 -113 1381
rect -45 1347 -29 1381
rect 29 1347 45 1381
rect 113 1347 129 1381
rect 187 1347 203 1381
rect 271 1347 287 1381
rect 345 1347 361 1381
rect 429 1347 445 1381
rect 503 1347 519 1381
rect 587 1347 603 1381
rect 661 1347 677 1381
rect 745 1347 761 1381
rect 819 1347 835 1381
rect 903 1347 919 1381
rect 977 1347 993 1381
rect 1061 1347 1077 1381
rect 1135 1347 1151 1381
rect 1219 1347 1235 1381
rect 1293 1347 1309 1381
rect 1377 1347 1393 1381
rect 1451 1347 1467 1381
rect 1535 1347 1551 1381
rect -1597 1288 -1563 1304
rect -1597 -1304 -1563 -1288
rect -1439 1288 -1405 1304
rect -1439 -1304 -1405 -1288
rect -1281 1288 -1247 1304
rect -1281 -1304 -1247 -1288
rect -1123 1288 -1089 1304
rect -1123 -1304 -1089 -1288
rect -965 1288 -931 1304
rect -965 -1304 -931 -1288
rect -807 1288 -773 1304
rect -807 -1304 -773 -1288
rect -649 1288 -615 1304
rect -649 -1304 -615 -1288
rect -491 1288 -457 1304
rect -491 -1304 -457 -1288
rect -333 1288 -299 1304
rect -333 -1304 -299 -1288
rect -175 1288 -141 1304
rect -175 -1304 -141 -1288
rect -17 1288 17 1304
rect -17 -1304 17 -1288
rect 141 1288 175 1304
rect 141 -1304 175 -1288
rect 299 1288 333 1304
rect 299 -1304 333 -1288
rect 457 1288 491 1304
rect 457 -1304 491 -1288
rect 615 1288 649 1304
rect 615 -1304 649 -1288
rect 773 1288 807 1304
rect 773 -1304 807 -1288
rect 931 1288 965 1304
rect 931 -1304 965 -1288
rect 1089 1288 1123 1304
rect 1089 -1304 1123 -1288
rect 1247 1288 1281 1304
rect 1247 -1304 1281 -1288
rect 1405 1288 1439 1304
rect 1405 -1304 1439 -1288
rect 1563 1288 1597 1304
rect 1563 -1304 1597 -1288
rect -1551 -1381 -1535 -1347
rect -1467 -1381 -1451 -1347
rect -1393 -1381 -1377 -1347
rect -1309 -1381 -1293 -1347
rect -1235 -1381 -1219 -1347
rect -1151 -1381 -1135 -1347
rect -1077 -1381 -1061 -1347
rect -993 -1381 -977 -1347
rect -919 -1381 -903 -1347
rect -835 -1381 -819 -1347
rect -761 -1381 -745 -1347
rect -677 -1381 -661 -1347
rect -603 -1381 -587 -1347
rect -519 -1381 -503 -1347
rect -445 -1381 -429 -1347
rect -361 -1381 -345 -1347
rect -287 -1381 -271 -1347
rect -203 -1381 -187 -1347
rect -129 -1381 -113 -1347
rect -45 -1381 -29 -1347
rect 29 -1381 45 -1347
rect 113 -1381 129 -1347
rect 187 -1381 203 -1347
rect 271 -1381 287 -1347
rect 345 -1381 361 -1347
rect 429 -1381 445 -1347
rect 503 -1381 519 -1347
rect 587 -1381 603 -1347
rect 661 -1381 677 -1347
rect 745 -1381 761 -1347
rect 819 -1381 835 -1347
rect 903 -1381 919 -1347
rect 977 -1381 993 -1347
rect 1061 -1381 1077 -1347
rect 1135 -1381 1151 -1347
rect 1219 -1381 1235 -1347
rect 1293 -1381 1309 -1347
rect 1377 -1381 1393 -1347
rect 1451 -1381 1467 -1347
rect 1535 -1381 1551 -1347
rect -1731 -1485 -1697 -1423
rect 1697 -1485 1731 -1423
rect -1731 -1519 -1635 -1485
rect 1635 -1519 1731 -1485
<< viali >>
rect -1535 1347 -1467 1381
rect -1377 1347 -1309 1381
rect -1219 1347 -1151 1381
rect -1061 1347 -993 1381
rect -903 1347 -835 1381
rect -745 1347 -677 1381
rect -587 1347 -519 1381
rect -429 1347 -361 1381
rect -271 1347 -203 1381
rect -113 1347 -45 1381
rect 45 1347 113 1381
rect 203 1347 271 1381
rect 361 1347 429 1381
rect 519 1347 587 1381
rect 677 1347 745 1381
rect 835 1347 903 1381
rect 993 1347 1061 1381
rect 1151 1347 1219 1381
rect 1309 1347 1377 1381
rect 1467 1347 1535 1381
rect -1597 -1288 -1563 1288
rect -1439 -1288 -1405 1288
rect -1281 -1288 -1247 1288
rect -1123 -1288 -1089 1288
rect -965 -1288 -931 1288
rect -807 -1288 -773 1288
rect -649 -1288 -615 1288
rect -491 -1288 -457 1288
rect -333 -1288 -299 1288
rect -175 -1288 -141 1288
rect -17 -1288 17 1288
rect 141 -1288 175 1288
rect 299 -1288 333 1288
rect 457 -1288 491 1288
rect 615 -1288 649 1288
rect 773 -1288 807 1288
rect 931 -1288 965 1288
rect 1089 -1288 1123 1288
rect 1247 -1288 1281 1288
rect 1405 -1288 1439 1288
rect 1563 -1288 1597 1288
rect -1535 -1381 -1467 -1347
rect -1377 -1381 -1309 -1347
rect -1219 -1381 -1151 -1347
rect -1061 -1381 -993 -1347
rect -903 -1381 -835 -1347
rect -745 -1381 -677 -1347
rect -587 -1381 -519 -1347
rect -429 -1381 -361 -1347
rect -271 -1381 -203 -1347
rect -113 -1381 -45 -1347
rect 45 -1381 113 -1347
rect 203 -1381 271 -1347
rect 361 -1381 429 -1347
rect 519 -1381 587 -1347
rect 677 -1381 745 -1347
rect 835 -1381 903 -1347
rect 993 -1381 1061 -1347
rect 1151 -1381 1219 -1347
rect 1309 -1381 1377 -1347
rect 1467 -1381 1535 -1347
<< metal1 >>
rect -1547 1381 -1455 1387
rect -1547 1347 -1535 1381
rect -1467 1347 -1455 1381
rect -1547 1341 -1455 1347
rect -1389 1381 -1297 1387
rect -1389 1347 -1377 1381
rect -1309 1347 -1297 1381
rect -1389 1341 -1297 1347
rect -1231 1381 -1139 1387
rect -1231 1347 -1219 1381
rect -1151 1347 -1139 1381
rect -1231 1341 -1139 1347
rect -1073 1381 -981 1387
rect -1073 1347 -1061 1381
rect -993 1347 -981 1381
rect -1073 1341 -981 1347
rect -915 1381 -823 1387
rect -915 1347 -903 1381
rect -835 1347 -823 1381
rect -915 1341 -823 1347
rect -757 1381 -665 1387
rect -757 1347 -745 1381
rect -677 1347 -665 1381
rect -757 1341 -665 1347
rect -599 1381 -507 1387
rect -599 1347 -587 1381
rect -519 1347 -507 1381
rect -599 1341 -507 1347
rect -441 1381 -349 1387
rect -441 1347 -429 1381
rect -361 1347 -349 1381
rect -441 1341 -349 1347
rect -283 1381 -191 1387
rect -283 1347 -271 1381
rect -203 1347 -191 1381
rect -283 1341 -191 1347
rect -125 1381 -33 1387
rect -125 1347 -113 1381
rect -45 1347 -33 1381
rect -125 1341 -33 1347
rect 33 1381 125 1387
rect 33 1347 45 1381
rect 113 1347 125 1381
rect 33 1341 125 1347
rect 191 1381 283 1387
rect 191 1347 203 1381
rect 271 1347 283 1381
rect 191 1341 283 1347
rect 349 1381 441 1387
rect 349 1347 361 1381
rect 429 1347 441 1381
rect 349 1341 441 1347
rect 507 1381 599 1387
rect 507 1347 519 1381
rect 587 1347 599 1381
rect 507 1341 599 1347
rect 665 1381 757 1387
rect 665 1347 677 1381
rect 745 1347 757 1381
rect 665 1341 757 1347
rect 823 1381 915 1387
rect 823 1347 835 1381
rect 903 1347 915 1381
rect 823 1341 915 1347
rect 981 1381 1073 1387
rect 981 1347 993 1381
rect 1061 1347 1073 1381
rect 981 1341 1073 1347
rect 1139 1381 1231 1387
rect 1139 1347 1151 1381
rect 1219 1347 1231 1381
rect 1139 1341 1231 1347
rect 1297 1381 1389 1387
rect 1297 1347 1309 1381
rect 1377 1347 1389 1381
rect 1297 1341 1389 1347
rect 1455 1381 1547 1387
rect 1455 1347 1467 1381
rect 1535 1347 1547 1381
rect 1455 1341 1547 1347
rect -1603 1288 -1557 1300
rect -1603 -1288 -1597 1288
rect -1563 -1288 -1557 1288
rect -1603 -1300 -1557 -1288
rect -1445 1288 -1399 1300
rect -1445 -1288 -1439 1288
rect -1405 -1288 -1399 1288
rect -1445 -1300 -1399 -1288
rect -1287 1288 -1241 1300
rect -1287 -1288 -1281 1288
rect -1247 -1288 -1241 1288
rect -1287 -1300 -1241 -1288
rect -1129 1288 -1083 1300
rect -1129 -1288 -1123 1288
rect -1089 -1288 -1083 1288
rect -1129 -1300 -1083 -1288
rect -971 1288 -925 1300
rect -971 -1288 -965 1288
rect -931 -1288 -925 1288
rect -971 -1300 -925 -1288
rect -813 1288 -767 1300
rect -813 -1288 -807 1288
rect -773 -1288 -767 1288
rect -813 -1300 -767 -1288
rect -655 1288 -609 1300
rect -655 -1288 -649 1288
rect -615 -1288 -609 1288
rect -655 -1300 -609 -1288
rect -497 1288 -451 1300
rect -497 -1288 -491 1288
rect -457 -1288 -451 1288
rect -497 -1300 -451 -1288
rect -339 1288 -293 1300
rect -339 -1288 -333 1288
rect -299 -1288 -293 1288
rect -339 -1300 -293 -1288
rect -181 1288 -135 1300
rect -181 -1288 -175 1288
rect -141 -1288 -135 1288
rect -181 -1300 -135 -1288
rect -23 1288 23 1300
rect -23 -1288 -17 1288
rect 17 -1288 23 1288
rect -23 -1300 23 -1288
rect 135 1288 181 1300
rect 135 -1288 141 1288
rect 175 -1288 181 1288
rect 135 -1300 181 -1288
rect 293 1288 339 1300
rect 293 -1288 299 1288
rect 333 -1288 339 1288
rect 293 -1300 339 -1288
rect 451 1288 497 1300
rect 451 -1288 457 1288
rect 491 -1288 497 1288
rect 451 -1300 497 -1288
rect 609 1288 655 1300
rect 609 -1288 615 1288
rect 649 -1288 655 1288
rect 609 -1300 655 -1288
rect 767 1288 813 1300
rect 767 -1288 773 1288
rect 807 -1288 813 1288
rect 767 -1300 813 -1288
rect 925 1288 971 1300
rect 925 -1288 931 1288
rect 965 -1288 971 1288
rect 925 -1300 971 -1288
rect 1083 1288 1129 1300
rect 1083 -1288 1089 1288
rect 1123 -1288 1129 1288
rect 1083 -1300 1129 -1288
rect 1241 1288 1287 1300
rect 1241 -1288 1247 1288
rect 1281 -1288 1287 1288
rect 1241 -1300 1287 -1288
rect 1399 1288 1445 1300
rect 1399 -1288 1405 1288
rect 1439 -1288 1445 1288
rect 1399 -1300 1445 -1288
rect 1557 1288 1603 1300
rect 1557 -1288 1563 1288
rect 1597 -1288 1603 1288
rect 1557 -1300 1603 -1288
rect -1547 -1347 -1455 -1341
rect -1547 -1381 -1535 -1347
rect -1467 -1381 -1455 -1347
rect -1547 -1387 -1455 -1381
rect -1389 -1347 -1297 -1341
rect -1389 -1381 -1377 -1347
rect -1309 -1381 -1297 -1347
rect -1389 -1387 -1297 -1381
rect -1231 -1347 -1139 -1341
rect -1231 -1381 -1219 -1347
rect -1151 -1381 -1139 -1347
rect -1231 -1387 -1139 -1381
rect -1073 -1347 -981 -1341
rect -1073 -1381 -1061 -1347
rect -993 -1381 -981 -1347
rect -1073 -1387 -981 -1381
rect -915 -1347 -823 -1341
rect -915 -1381 -903 -1347
rect -835 -1381 -823 -1347
rect -915 -1387 -823 -1381
rect -757 -1347 -665 -1341
rect -757 -1381 -745 -1347
rect -677 -1381 -665 -1347
rect -757 -1387 -665 -1381
rect -599 -1347 -507 -1341
rect -599 -1381 -587 -1347
rect -519 -1381 -507 -1347
rect -599 -1387 -507 -1381
rect -441 -1347 -349 -1341
rect -441 -1381 -429 -1347
rect -361 -1381 -349 -1347
rect -441 -1387 -349 -1381
rect -283 -1347 -191 -1341
rect -283 -1381 -271 -1347
rect -203 -1381 -191 -1347
rect -283 -1387 -191 -1381
rect -125 -1347 -33 -1341
rect -125 -1381 -113 -1347
rect -45 -1381 -33 -1347
rect -125 -1387 -33 -1381
rect 33 -1347 125 -1341
rect 33 -1381 45 -1347
rect 113 -1381 125 -1347
rect 33 -1387 125 -1381
rect 191 -1347 283 -1341
rect 191 -1381 203 -1347
rect 271 -1381 283 -1347
rect 191 -1387 283 -1381
rect 349 -1347 441 -1341
rect 349 -1381 361 -1347
rect 429 -1381 441 -1347
rect 349 -1387 441 -1381
rect 507 -1347 599 -1341
rect 507 -1381 519 -1347
rect 587 -1381 599 -1347
rect 507 -1387 599 -1381
rect 665 -1347 757 -1341
rect 665 -1381 677 -1347
rect 745 -1381 757 -1347
rect 665 -1387 757 -1381
rect 823 -1347 915 -1341
rect 823 -1381 835 -1347
rect 903 -1381 915 -1347
rect 823 -1387 915 -1381
rect 981 -1347 1073 -1341
rect 981 -1381 993 -1347
rect 1061 -1381 1073 -1347
rect 981 -1387 1073 -1381
rect 1139 -1347 1231 -1341
rect 1139 -1381 1151 -1347
rect 1219 -1381 1231 -1347
rect 1139 -1387 1231 -1381
rect 1297 -1347 1389 -1341
rect 1297 -1381 1309 -1347
rect 1377 -1381 1389 -1347
rect 1297 -1387 1389 -1381
rect 1455 -1347 1547 -1341
rect 1455 -1381 1467 -1347
rect 1535 -1381 1547 -1347
rect 1455 -1387 1547 -1381
<< properties >>
string FIXED_BBOX -1714 -1502 1714 1502
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 13.0 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
