magic
tech sky130A
magscale 1 2
timestamp 1697185551
<< viali >>
rect 1324 2182 1358 2556
rect 128 1590 370 1624
<< metal1 >>
rect -66 3062 1228 3492
rect -68 2552 456 2620
rect -68 2248 102 2552
rect 280 2248 456 2552
rect -68 2190 456 2248
rect 704 2570 1228 2622
rect 704 2266 880 2570
rect 1058 2266 1228 2570
rect 704 2192 1228 2266
rect 1312 2556 1566 2568
rect 1312 2182 1324 2556
rect 1358 2182 1566 2556
rect 1312 2170 1566 2182
rect 116 1634 382 1638
rect 116 1582 126 1634
rect 376 1582 382 1634
rect 116 1578 382 1582
rect 1394 1498 1568 2170
rect 84 1468 1664 1498
rect 84 1456 286 1468
rect 84 1220 286 1234
rect 320 1220 354 1468
rect 507 1456 720 1468
rect 507 1450 707 1456
rect 754 1440 788 1468
rect 945 1456 1158 1468
rect 945 1450 1145 1456
rect 1192 1440 1226 1468
rect 1383 1456 1596 1468
rect 1383 1450 1583 1456
rect 1630 1440 1664 1468
rect 748 1248 794 1440
rect 1186 1248 1232 1440
rect 1624 1248 1670 1440
rect 84 1192 354 1220
rect 507 1234 707 1238
rect 507 1220 720 1234
rect 754 1220 788 1248
rect 507 1192 788 1220
rect 945 1234 1145 1238
rect 945 1220 1158 1234
rect 1192 1220 1226 1248
rect 945 1192 1226 1220
rect 1383 1234 1583 1238
rect 1383 1220 1596 1234
rect 1630 1220 1664 1248
rect 1383 1192 1664 1220
rect 320 1120 354 1192
rect 84 1118 354 1120
rect 73 1090 354 1118
rect 73 1078 286 1090
rect 73 1072 273 1078
rect 320 1062 354 1090
rect 508 1130 710 1136
rect 508 1072 514 1130
rect 704 1072 710 1130
rect 508 1066 710 1072
rect 944 1130 1146 1136
rect 944 1072 950 1130
rect 1140 1072 1146 1130
rect 1628 1120 1664 1192
rect 1392 1118 1664 1120
rect 1381 1090 1664 1118
rect 1381 1078 1594 1090
rect 1381 1072 1581 1078
rect 944 1066 1146 1072
rect 1628 1066 1664 1090
rect 1628 1062 1668 1066
rect 314 870 360 1062
rect 502 902 710 908
rect 73 856 273 860
rect 73 842 286 856
rect 320 842 354 870
rect 73 814 354 842
rect 502 814 508 902
rect 704 860 710 902
rect 750 880 904 1062
rect 738 870 904 880
rect 1622 870 1668 1062
rect 738 860 852 870
rect 704 814 852 860
rect 320 742 354 814
rect 508 808 710 814
rect 84 740 354 742
rect 932 740 1146 862
rect 1381 856 1581 860
rect 1381 842 1594 856
rect 1628 842 1664 870
rect 1381 814 1664 842
rect 1630 740 1664 814
rect 73 712 354 740
rect 709 738 1146 740
rect 73 700 286 712
rect 73 694 273 700
rect 320 680 354 712
rect 510 712 1146 738
rect 510 694 722 712
rect 932 692 1146 712
rect 1392 712 1664 740
rect 1392 700 1594 712
rect 1630 684 1664 712
rect 314 492 360 680
rect 416 678 480 684
rect 416 498 422 678
rect 1178 676 1250 678
rect 416 492 480 498
rect 508 494 710 500
rect 320 488 354 492
rect 73 478 273 482
rect 73 464 286 478
rect 320 464 352 488
rect 73 436 352 464
rect 318 364 352 436
rect 508 436 514 494
rect 704 436 710 494
rect 508 430 710 436
rect 944 494 1146 500
rect 1178 496 1186 676
rect 1244 496 1250 676
rect 1178 494 1250 496
rect 944 436 950 494
rect 1140 478 1146 494
rect 1628 492 1664 684
rect 1140 436 1150 478
rect 1392 464 1594 476
rect 1630 464 1664 492
rect 1392 436 1664 464
rect 944 430 1146 436
rect 1630 364 1664 436
rect 82 362 352 364
rect 520 362 790 364
rect 954 362 1224 364
rect 1394 362 1664 364
rect 71 334 352 362
rect 71 322 284 334
rect 71 316 271 322
rect 318 306 352 334
rect 509 334 790 362
rect 509 322 722 334
rect 509 316 709 322
rect 756 306 790 334
rect 943 334 1224 362
rect 943 322 1156 334
rect 943 316 1143 322
rect 1190 306 1224 334
rect 1383 334 1664 362
rect 1383 322 1596 334
rect 1383 316 1583 322
rect 1630 306 1664 334
rect 312 114 358 306
rect 750 114 796 306
rect 1184 114 1230 306
rect 1624 114 1670 306
rect 71 100 271 104
rect 71 86 284 100
rect 318 86 352 114
rect 509 100 709 104
rect 506 86 722 100
rect 756 86 790 114
rect 943 100 1143 104
rect 943 86 1156 100
rect 1190 86 1224 114
rect 1368 86 1594 104
rect 1630 86 1664 114
rect 71 58 1664 86
<< via1 >>
rect 102 2248 280 2552
rect 880 2266 1058 2570
rect 126 1624 376 1634
rect 126 1590 128 1624
rect 128 1590 370 1624
rect 370 1590 376 1624
rect 126 1582 376 1590
rect 514 1072 704 1130
rect 950 1072 1140 1130
rect 508 814 704 902
rect 422 498 480 678
rect 514 436 704 494
rect 1186 496 1244 676
rect 950 436 1140 494
<< metal2 >>
rect 874 2574 1066 2576
rect 874 2570 1146 2574
rect 92 2552 292 2560
rect 92 2248 102 2552
rect 280 2248 292 2552
rect 874 2266 880 2570
rect 1058 2266 1146 2570
rect 874 2258 1146 2266
rect 92 1934 292 2248
rect -490 1924 292 1934
rect -490 1776 710 1924
rect 944 1892 1146 2258
rect 944 1880 1148 1892
rect 508 1638 710 1776
rect 120 1634 710 1638
rect 120 1582 126 1634
rect 376 1582 710 1634
rect 120 1578 710 1582
rect 508 1130 710 1578
rect 946 1136 1148 1880
rect 508 1072 514 1130
rect 704 1072 710 1130
rect 508 1064 710 1072
rect 944 1130 1148 1136
rect 944 1072 950 1130
rect 1140 1072 1148 1130
rect 944 1068 1148 1072
rect 944 1066 1146 1068
rect -444 902 712 918
rect -444 814 508 902
rect 704 814 712 902
rect -444 806 712 814
rect 416 680 480 684
rect -430 678 480 680
rect -430 498 422 678
rect 1178 680 1998 682
rect 1178 676 2222 680
rect -430 492 480 498
rect 508 500 708 504
rect 508 494 710 500
rect 944 498 1146 500
rect 508 470 514 494
rect 506 436 514 470
rect 704 436 710 494
rect 506 430 710 436
rect 942 494 1146 498
rect 1178 496 1186 676
rect 1244 496 2222 676
rect 1178 494 2222 496
rect 942 436 950 494
rect 1140 436 1146 494
rect 1700 492 1810 494
rect 942 430 1146 436
rect 506 -508 708 430
rect 942 -514 1144 430
use sky130_fd_pr__pfet_g5v0d10v5_XGMD62  sky130_fd_pr__pfet_g5v0d10v5_XGMD62_0
timestamp 1696881349
transform 0 -1 827 1 0 777
box -925 -1051 925 1051
use sky130_fd_pr__res_xhigh_po_0p69_XDW3D2#0  sky130_fd_pr__res_xhigh_po_0p69_XDW3D2_0
timestamp 1696354057
transform 1 0 581 0 1 2841
box -814 -818 814 818
<< labels >>
rlabel metal2 -462 1800 -102 1908 1 vsup
port 1 n
rlabel metal2 554 -468 648 -254 1 iout
port 4 n
rlabel metal2 998 -470 1092 -256 1 iout_n
port 5 n
rlabel metal2 1832 546 2064 640 1 vbias
port 7 n
rlabel metal2 -422 816 -156 908 1 iref
port 3 n
rlabel metal2 -368 538 -136 632 1 vsw
port 6 n
rlabel metal1 1378 2216 1536 2530 3 vgnd
<< end >>
