magic
tech sky130A
magscale 1 2
timestamp 1628516087
<< metal1 >>
rect 16 4694 7368 5694
rect 192 3904 242 4694
rect 774 4368 830 4694
rect 2006 4396 2062 4694
rect 646 4366 990 4368
rect 646 4314 989 4366
rect 1041 4314 1047 4366
rect 1832 4340 2175 4396
rect 2227 4342 2233 4394
rect 646 4312 990 4314
rect 646 4150 702 4312
rect 1832 4178 1888 4340
rect 2174 4160 2226 4166
rect 988 4132 1040 4138
rect 2174 4102 2226 4108
rect 988 4074 1040 4080
rect 990 4000 1037 4074
rect 2176 4028 2223 4102
rect -1226 3146 -883 3202
rect -831 3148 -825 3200
rect -1226 2984 -1170 3146
rect -884 2966 -832 2972
rect -884 2908 -832 2914
rect 832 2910 879 2984
rect 2018 2912 2065 2986
rect -882 2834 -835 2908
rect 829 2904 881 2910
rect 829 2846 881 2852
rect 2015 2906 2067 2912
rect 2015 2848 2067 2854
rect 1167 2756 1223 2834
rect 730 2710 2324 2756
rect 1167 2672 1223 2710
rect 2353 2674 2409 2836
rect 822 2618 828 2670
rect 880 2616 1223 2672
rect 2008 2620 2014 2672
rect 2066 2618 2409 2674
rect 970 2398 1026 2616
rect 2202 2398 2258 2618
rect 712 2342 1026 2398
rect 1472 2342 2258 2398
rect 432 2180 552 2252
rect 624 2180 630 2252
rect 432 1706 504 2180
rect 712 1878 768 2342
rect 216 1634 504 1706
rect 898 908 1342 1908
rect 1472 1878 1528 2342
rect 1908 2124 2000 2130
rect 1908 1940 2000 2032
rect 2466 2014 2658 2020
rect 2466 1942 2586 2014
rect 2466 1940 2658 1942
rect 796 336 888 830
rect 1084 484 1156 908
rect 1084 406 1156 412
rect 54 -64 888 336
rect 1352 -92 1444 830
rect 1664 134 1670 206
rect 1742 134 1886 206
rect 2010 -92 2456 1908
rect 2586 1836 2658 1940
rect 6275 1864 6281 1941
rect 6358 1864 6364 1941
rect 6281 1670 6358 1864
rect 6281 1626 7174 1670
rect 6290 1624 7174 1626
rect 8398 301 8444 337
rect 8395 295 8447 301
rect 8395 237 8447 243
rect 6394 136 6440 172
rect 6711 138 6757 174
rect 7027 142 7073 178
rect 6391 130 6443 136
rect 6391 72 6443 78
rect 6708 132 6760 138
rect 6708 74 6760 80
rect 7024 136 7076 142
rect 7024 78 7076 84
rect 54 -492 1444 -92
rect 2197 -548 2269 -92
rect 6704 -190 6710 -138
rect 6762 -190 6768 -138
rect 6713 -548 6759 -190
rect 54 -1548 7406 -548
<< via1 >>
rect 989 4314 1041 4366
rect 2175 4342 2227 4394
rect 988 4080 1040 4132
rect 2174 4108 2226 4160
rect -883 3148 -831 3200
rect -884 2914 -832 2966
rect 829 2852 881 2904
rect 2015 2854 2067 2906
rect 828 2618 880 2670
rect 2014 2620 2066 2672
rect 552 2180 624 2252
rect 1908 2032 2000 2124
rect 2586 1942 2658 2014
rect 1084 412 1156 484
rect 1670 134 1742 206
rect 6281 1864 6358 1941
rect 8395 243 8447 295
rect 6391 78 6443 130
rect 6708 80 6760 132
rect 7024 84 7076 136
rect 6710 -190 6762 -138
<< metal2 >>
rect 2175 4394 2227 4400
rect 989 4366 1041 4372
rect 2175 4336 2227 4342
rect 989 4308 1041 4314
rect 991 4132 1038 4308
rect 2177 4160 2224 4336
rect 982 4080 988 4132
rect 1040 4080 1046 4132
rect 2168 4108 2174 4160
rect 2226 4108 2232 4160
rect -883 3200 -831 3206
rect -883 3142 -831 3148
rect -881 2966 -834 3142
rect -890 2914 -884 2966
rect -832 2914 -826 2966
rect 823 2852 829 2904
rect 881 2852 887 2904
rect 2009 2854 2015 2906
rect 2067 2854 2073 2906
rect 831 2676 878 2852
rect 2017 2678 2064 2854
rect 828 2670 880 2676
rect 828 2612 880 2618
rect 2014 2672 2066 2678
rect 2014 2614 2066 2620
rect 552 2252 624 2258
rect 624 2180 2658 2252
rect 552 2174 624 2180
rect 1908 2124 2000 2180
rect 1902 2032 1908 2124
rect 2000 2032 2006 2124
rect 2586 2019 2658 2180
rect 2586 2014 2838 2019
rect 2580 1942 2586 2014
rect 2658 1942 2838 2014
rect 2761 1941 2838 1942
rect 6281 1941 6358 1947
rect 2761 1864 6281 1941
rect 6281 1858 6358 1864
rect 1078 412 1084 484
rect 1156 412 1162 484
rect 1084 206 1156 412
rect 8389 243 8395 295
rect 8447 243 8453 295
rect 1670 206 1742 212
rect 1084 134 1670 206
rect 1670 128 1742 134
rect 6385 78 6391 130
rect 6443 78 6449 130
rect 6702 80 6708 132
rect 6760 80 6766 132
rect 7018 84 7024 136
rect 7076 84 7082 136
rect 6394 -141 6440 78
rect 6711 -132 6757 80
rect 6710 -138 6762 -132
rect 6394 -187 6710 -141
rect 7027 -141 7073 84
rect 8398 12 8444 243
rect 6762 -187 7073 -141
rect 6710 -196 6762 -190
use sky130_fd_pr__res_xhigh_po_0p35_X24WYH  sky130_fd_pr__res_xhigh_po_0p35_X24WYH_0
timestamp 1628260645
transform -1 0 217 0 1 2896
box -201 -1598 201 1598
use sky130_fd_pr__nfet_g5v0d10v5_A263FC  sky130_fd_pr__nfet_g5v0d10v5_A263FC_0
timestamp 1628499526
transform 1 0 842 0 1 1408
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_A263FC  sky130_fd_pr__nfet_g5v0d10v5_A263FC_1
timestamp 1628499526
transform 1 0 1398 0 1 1408
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_6HNVDQ  sky130_fd_pr__nfet_g5v0d10v5_6HNVDQ_0
timestamp 1628499526
transform 1 0 1954 0 1 908
box -278 -1258 278 1258
use sky130_fd_pr__nfet_g5v0d10v5_6HNVDQ  sky130_fd_pr__nfet_g5v0d10v5_6HNVDQ_1
timestamp 1628499526
transform 1 0 2512 0 1 908
box -278 -1258 278 1258
use sky130_fd_pr__cap_mim_m3_1_V36R79  sky130_fd_pr__cap_mim_m3_1_V36R79_0
timestamp 1628238145
transform 1 0 4460 0 1 750
box -1550 -1100 1549 1100
use sky130_fd_pr__pfet_g5v0d10v5_FGZEPY  sky130_fd_pr__pfet_g5v0d10v5_FGZEPY_0
timestamp 1628235263
transform 1 0 5123 0 1 3197
box -2283 -1297 2283 1297
use sky130_fd_pr__nfet_g5v0d10v5_USLVMX  sky130_fd_pr__nfet_g5v0d10v5_USLVMX_0
timestamp 1628499526
transform 1 0 6733 0 1 792
box -673 -1058 673 1058
use sky130_fd_pr__pfet_g5v0d10v5_WLXSDU  sky130_fd_pr__pfet_g5v0d10v5_WLXSDU_1
timestamp 1628235263
transform 1 0 934 0 1 3497
box -466 -997 466 997
use sky130_fd_pr__pfet_g5v0d10v5_WLXSDU  sky130_fd_pr__pfet_g5v0d10v5_WLXSDU_0
timestamp 1628235263
transform 1 0 2120 0 1 3497
box -466 -997 466 997
<< labels >>
rlabel metal1 54 -1548 7406 -548 0 ground
rlabel metal1 54 -492 984 -92 0 inNeg
rlabel space 54 -64 984 336 0 inPos
rlabel metal1 16 4694 7368 5694 0 power
<< end >>
