magic
tech sky130A
magscale 1 2
timestamp 1697652271
<< pwell >>
rect -739 -868 739 868
<< psubdiff >>
rect -703 798 -607 832
rect 607 798 703 832
rect -703 736 -669 798
rect 669 736 703 798
rect -703 -798 -669 -736
rect 669 -798 703 -736
rect -703 -832 -607 -798
rect 607 -832 703 -798
<< psubdiffcont >>
rect -607 798 607 832
rect -703 -736 -669 736
rect 669 -736 703 736
rect -607 -832 607 -798
<< xpolycontact >>
rect -573 270 573 702
rect -573 -702 573 -270
<< xpolyres >>
rect -573 -270 573 270
<< locali >>
rect -703 798 -607 832
rect 607 798 703 832
rect -703 736 -669 798
rect 669 736 703 798
rect -703 -798 -669 -736
rect 669 -798 703 -736
rect -703 -832 -607 -798
rect 607 -832 703 -798
<< viali >>
rect -557 287 557 684
rect -557 -684 557 -287
<< metal1 >>
rect -569 684 569 690
rect -569 287 -557 684
rect 557 287 569 684
rect -569 281 569 287
rect -569 -287 569 -281
rect -569 -684 -557 -287
rect 557 -684 569 -287
rect -569 -690 569 -684
<< res5p73 >>
rect -575 -272 575 272
<< properties >>
string FIXED_BBOX -686 -815 686 815
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 2.7 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 1.008k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
