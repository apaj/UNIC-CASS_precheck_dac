magic
tech sky130A
magscale 1 2
timestamp 1628235594
<< pwell >>
rect -278 -2585 278 2585
<< nnmos >>
rect -50 1327 50 2327
rect -50 109 50 1109
rect -50 -1109 50 -109
rect -50 -2327 50 -1327
<< mvndiff >>
rect -108 2315 -50 2327
rect -108 1339 -96 2315
rect -62 1339 -50 2315
rect -108 1327 -50 1339
rect 50 2315 108 2327
rect 50 1339 62 2315
rect 96 1339 108 2315
rect 50 1327 108 1339
rect -108 1097 -50 1109
rect -108 121 -96 1097
rect -62 121 -50 1097
rect -108 109 -50 121
rect 50 1097 108 1109
rect 50 121 62 1097
rect 96 121 108 1097
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -1097 -96 -121
rect -62 -1097 -50 -121
rect -108 -1109 -50 -1097
rect 50 -121 108 -109
rect 50 -1097 62 -121
rect 96 -1097 108 -121
rect 50 -1109 108 -1097
rect -108 -1339 -50 -1327
rect -108 -2315 -96 -1339
rect -62 -2315 -50 -1339
rect -108 -2327 -50 -2315
rect 50 -1339 108 -1327
rect 50 -2315 62 -1339
rect 96 -2315 108 -1339
rect 50 -2327 108 -2315
<< mvndiffc >>
rect -96 1339 -62 2315
rect 62 1339 96 2315
rect -96 121 -62 1097
rect 62 121 96 1097
rect -96 -1097 -62 -121
rect 62 -1097 96 -121
rect -96 -2315 -62 -1339
rect 62 -2315 96 -1339
<< mvpsubdiff >>
rect -242 2537 242 2549
rect -242 2503 -134 2537
rect 134 2503 242 2537
rect -242 2491 242 2503
rect -242 2441 -184 2491
rect -242 -2441 -230 2441
rect -196 -2441 -184 2441
rect 184 2441 242 2491
rect -242 -2491 -184 -2441
rect 184 -2441 196 2441
rect 230 -2441 242 2441
rect 184 -2491 242 -2441
rect -242 -2503 242 -2491
rect -242 -2537 -134 -2503
rect 134 -2537 242 -2503
rect -242 -2549 242 -2537
<< mvpsubdiffcont >>
rect -134 2503 134 2537
rect -230 -2441 -196 2441
rect 196 -2441 230 2441
rect -134 -2537 134 -2503
<< poly >>
rect -50 2399 50 2415
rect -50 2365 -34 2399
rect 34 2365 50 2399
rect -50 2327 50 2365
rect -50 1289 50 1327
rect -50 1255 -34 1289
rect 34 1255 50 1289
rect -50 1239 50 1255
rect -50 1181 50 1197
rect -50 1147 -34 1181
rect 34 1147 50 1181
rect -50 1109 50 1147
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -1147 50 -1109
rect -50 -1181 -34 -1147
rect 34 -1181 50 -1147
rect -50 -1197 50 -1181
rect -50 -1255 50 -1239
rect -50 -1289 -34 -1255
rect 34 -1289 50 -1255
rect -50 -1327 50 -1289
rect -50 -2365 50 -2327
rect -50 -2399 -34 -2365
rect 34 -2399 50 -2365
rect -50 -2415 50 -2399
<< polycont >>
rect -34 2365 34 2399
rect -34 1255 34 1289
rect -34 1147 34 1181
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -1181 34 -1147
rect -34 -1289 34 -1255
rect -34 -2399 34 -2365
<< locali >>
rect -230 2503 -134 2537
rect 134 2503 230 2537
rect -230 2441 -196 2503
rect 196 2441 230 2503
rect -50 2365 -34 2399
rect 34 2365 50 2399
rect -96 2315 -62 2331
rect -96 1323 -62 1339
rect 62 2315 96 2331
rect 62 1323 96 1339
rect -50 1255 -34 1289
rect 34 1255 50 1289
rect -50 1147 -34 1181
rect 34 1147 50 1181
rect -96 1097 -62 1113
rect -96 105 -62 121
rect 62 1097 96 1113
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -1113 -62 -1097
rect 62 -121 96 -105
rect 62 -1113 96 -1097
rect -50 -1181 -34 -1147
rect 34 -1181 50 -1147
rect -50 -1289 -34 -1255
rect 34 -1289 50 -1255
rect -96 -1339 -62 -1323
rect -96 -2331 -62 -2315
rect 62 -1339 96 -1323
rect 62 -2331 96 -2315
rect -50 -2399 -34 -2365
rect 34 -2399 50 -2365
rect -230 -2503 -196 -2441
rect 196 -2503 230 -2441
rect -230 -2537 -134 -2503
rect 134 -2537 230 -2503
<< viali >>
rect -34 2365 34 2399
rect -96 1339 -62 2315
rect 62 1339 96 2315
rect -34 1255 34 1289
rect -34 1147 34 1181
rect -96 121 -62 1097
rect 62 121 96 1097
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -1097 -62 -121
rect 62 -1097 96 -121
rect -34 -1181 34 -1147
rect -34 -1289 34 -1255
rect -96 -2315 -62 -1339
rect 62 -2315 96 -1339
rect -34 -2399 34 -2365
<< metal1 >>
rect -46 2399 46 2405
rect -46 2365 -34 2399
rect 34 2365 46 2399
rect -46 2359 46 2365
rect -102 2315 -56 2327
rect -102 1339 -96 2315
rect -62 1339 -56 2315
rect -102 1327 -56 1339
rect 56 2315 102 2327
rect 56 1339 62 2315
rect 96 1339 102 2315
rect 56 1327 102 1339
rect -46 1289 46 1295
rect -46 1255 -34 1289
rect 34 1255 46 1289
rect -46 1249 46 1255
rect -46 1181 46 1187
rect -46 1147 -34 1181
rect 34 1147 46 1181
rect -46 1141 46 1147
rect -102 1097 -56 1109
rect -102 121 -96 1097
rect -62 121 -56 1097
rect -102 109 -56 121
rect 56 1097 102 1109
rect 56 121 62 1097
rect 96 121 102 1097
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -1097 -96 -121
rect -62 -1097 -56 -121
rect -102 -1109 -56 -1097
rect 56 -121 102 -109
rect 56 -1097 62 -121
rect 96 -1097 102 -121
rect 56 -1109 102 -1097
rect -46 -1147 46 -1141
rect -46 -1181 -34 -1147
rect 34 -1181 46 -1147
rect -46 -1187 46 -1181
rect -46 -1255 46 -1249
rect -46 -1289 -34 -1255
rect 34 -1289 46 -1255
rect -46 -1295 46 -1289
rect -102 -1339 -56 -1327
rect -102 -2315 -96 -1339
rect -62 -2315 -56 -1339
rect -102 -2327 -56 -2315
rect 56 -1339 102 -1327
rect 56 -2315 62 -1339
rect 96 -2315 102 -1339
rect 56 -2327 102 -2315
rect -46 -2365 46 -2359
rect -46 -2399 -34 -2365
rect 34 -2399 46 -2365
rect -46 -2405 46 -2399
<< properties >>
string gencell sky130_fd_pr__nfet_03v3_nvt
string FIXED_BBOX -213 -2520 213 2520
string parameters w 5 l 0.50 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
