magic
tech sky130A
magscale 1 2
timestamp 1628238145
<< metal3 >>
rect -1550 1072 1549 1100
rect -1550 -1072 1465 1072
rect 1529 -1072 1549 1072
rect -1550 -1100 1549 -1072
<< via3 >>
rect 1465 -1072 1529 1072
<< mimcap >>
rect -1450 960 1350 1000
rect -1450 -960 -1410 960
rect 1310 -960 1350 960
rect -1450 -1000 1350 -960
<< mimcapcontact >>
rect -1410 -960 1310 960
<< metal4 >>
rect 1449 1072 1545 1088
rect -1411 960 1311 961
rect -1411 -960 -1410 960
rect 1310 -960 1311 960
rect -1411 -961 1311 -960
rect 1449 -1072 1465 1072
rect 1529 -1072 1545 1072
rect 1449 -1088 1545 -1072
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -1550 -1100 1450 1100
string parameters w 14 l 10 val 289.12 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
