* NGSPICE file created from dac_top_cell.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p69_RV3JGD a_n69_1300# a_n69_n1732# a_n199_n1862#
X0 a_n69_n1732# a_n69_1300# a_n199_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGUWVM a_n100_n197# a_100_n100# w_n358_n397#
+ a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n358_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGR8VM a_n100_n497# a_100_n400# w_n358_n697#
+ a_n158_n400#
X0 a_100_n400# a_n100_n497# a_n158_n400# w_n358_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt dac_cell3 vsup iref vsw iout iout_n vbias vgnd
XXR1 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69_RV3JGD
XXR2 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69_RV3JGD
XXR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69_RV3JGD
XXR4 vsup parR vgnd sky130_fd_pr__res_xhigh_po_0p69_RV3JGD
XXM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5_FGUWVM
XXM2 iref sourceM3M4 vsup sourceM2 sky130_fd_pr__pfet_g5v0d10v5_FGR8VM
XXM3 vsw iout vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGR8VM
XXM4 vbias iout_n vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGR8VM
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_MS44J6 a_n69_n6232# a_n69_5800# a_n199_n6362#
X0 a_n69_n6232# a_n69_5800# a_n199_n6362# sky130_fd_pr__res_xhigh_po_0p69 l=58
.ends

.subckt dac_cell1 vsup iref vsw iout iout_n vbias vgnd
XXR1 parR sourceM2 vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXR2 parR sourceM2 vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXR4 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5_FGUWVM
XXM2 iref sourceM3M4 vsup sourceM2 sky130_fd_pr__pfet_g5v0d10v5_FGUWVM
XXM3 vsw iout vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGUWVM
XXM4 vbias iout_n vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGUWVM
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_5CVACY a_n199_n1162# a_n69_600# a_n69_n1032#
X0 a_n69_600# a_n69_n1032# a_n199_n1162# sky130_fd_pr__res_xhigh_po_0p69 l=6
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y a_50_n500# a_n242_n722# a_n108_n500# a_n50_n588#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n242_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NQCFE9 a_189_n500# a_89_n588# a_31_n500# a_n189_n588#
+ a_n381_n722# a_n89_n500# a_n247_n500#
X0 a_189_n500# a_89_n588# a_31_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
X1 a_n89_n500# a_n189_n588# a_n247_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CJGAEC a_189_n500# a_89_n588# a_31_n500# a_n189_n588#
+ a_n381_n722# a_n89_n500# a_n247_n500#
X0 a_189_n500# a_89_n588# a_31_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
X1 a_n89_n500# a_n189_n588# a_n247_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2MGL8M a_367_n688# a_89_n688# a_31_n600# a_n189_n688#
+ a_n1023_n688# a_645_n688# a_n467_n688# a_923_n688# a_n745_n688# a_n89_n600# a_n367_n600#
+ a_n645_n600# a_n1081_n600# a_n247_n600# a_n923_n600# a_n525_n600# a_n803_n600# a_309_n600#
+ a_587_n600# a_189_n600# a_865_n600# a_467_n600# a_n1215_n822# a_745_n600# a_1023_n600#
X0 a_n367_n600# a_n467_n688# a_n525_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X1 a_467_n600# a_367_n688# a_309_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X2 a_189_n600# a_89_n688# a_31_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X3 a_n645_n600# a_n745_n688# a_n803_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X4 a_745_n600# a_645_n688# a_587_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X5 a_n89_n600# a_n189_n688# a_n247_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X6 a_n923_n600# a_n1023_n688# a_n1081_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X7 a_1023_n600# a_923_n688# a_865_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_X3UTN5 a_170_n700# a_n50_n797# a_50_n700# a_n228_n700#
+ w_n586_n997# a_n108_n700# a_n386_n700# a_228_n797# a_n328_n797# a_328_n700#
X0 a_328_n700# a_228_n797# a_170_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X1 a_50_n700# a_n50_n797# a_n108_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X2 a_n228_n700# a_n328_n797# a_n386_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AE43MT a_170_n700# a_n50_n797# a_50_n700# a_n228_n700#
+ w_n586_n997# a_n108_n700# a_n386_n700# a_228_n797# a_n328_n797# a_328_n700#
X0 a_328_n700# a_228_n797# a_170_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X1 a_50_n700# a_n50_n797# a_n108_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X2 a_n228_n700# a_n328_n797# a_n386_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CNRWF7 a_1579_n1300# a_n803_n1300# a_n1757_n1300#
+ a_n2035_n1300# a_1301_n1300# a_n645_n1300# a_1143_n1300# a_n2413_n1397# a_n2691_n1397#
+ a_n1637_n1300# a_n2193_n1300# a_189_n1300# a_n525_n1300# a_2591_n1397# a_2313_n1397#
+ a_923_n1397# a_2533_n1300# a_1023_n1300# a_n1479_n1300# a_n367_n1300# a_n1201_n1300#
+ a_n1857_n1397# a_n2135_n1397# a_n745_n1397# a_2691_n1300# a_2413_n1300# a_n89_n1300#
+ a_n1359_n1300# a_n247_n1300# a_645_n1397# a_2255_n1300# a_1977_n1300# a_865_n1300#
+ a_2035_n1397# a_1757_n1397# a_n2749_n1300# a_n1579_n1397# a_n1301_n1397# a_2135_n1300#
+ a_1857_n1300# a_745_n1300# a_n467_n1397# a_n1081_n1300# a_n2313_n1300# a_n2591_n1300#
+ a_89_n1397# a_587_n1300# a_309_n1300# a_1479_n1397# a_367_n1397# a_1699_n1300# a_31_n1300#
+ a_n923_n1300# a_1201_n1397# a_1421_n1300# a_n1915_n1300# a_n2471_n1300# a_467_n1300#
+ a_n189_n1397# a_n1023_n1397#
X0 a_1857_n1300# a_1757_n1397# a_1699_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X1 a_2691_n1300# a_2591_n1397# a_2533_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X2 a_n923_n1300# a_n1023_n1397# a_n1081_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X3 a_745_n1300# a_645_n1397# a_587_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X4 a_n2035_n1300# a_n2135_n1397# a_n2193_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X5 a_1579_n1300# a_1479_n1397# a_1421_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X6 a_467_n1300# a_367_n1397# a_309_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X7 a_n645_n1300# a_n745_n1397# a_n803_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X8 a_n2591_n1300# a_n2691_n1397# a_n2749_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X9 a_n1757_n1300# a_n1857_n1397# a_n1915_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X10 a_n367_n1300# a_n467_n1397# a_n525_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X11 a_1301_n1300# a_1201_n1397# a_1143_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X12 a_2413_n1300# a_2313_n1397# a_2255_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X13 a_n1479_n1300# a_n1579_n1397# a_n1637_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X14 a_n89_n1300# a_n189_n1397# a_n247_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X15 a_2135_n1300# a_2035_n1397# a_1977_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X16 a_189_n1300# a_89_n1397# a_31_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X17 a_n1201_n1300# a_n1301_n1397# a_n1359_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X18 a_1023_n1300# a_923_n1397# a_865_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X19 a_n2313_n1300# a_n2413_n1397# a_n2471_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_C5B489
X0 c1_n1050_n1400# m3_n1150_n1500# sky130_fd_pr__cap_mim_m3_1 l=14 w=10
.ends

.subckt miel21_opamp inPos inNeg outSingle power ground VSUBS
XXR1 VSUBS m1_n1838_8400# ground sky130_fd_pr__res_xhigh_po_0p69_5CVACY
XXR2 VSUBS m1_n1838_8400# m1_360_8394# sky130_fd_pr__res_xhigh_po_0p69_5CVACY
XXR3 VSUBS m1_360_8394# power sky130_fd_pr__res_xhigh_po_0p69_5CVACY
XXM1 m1_n536_4966# VSUBS ground inPos sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM2 m1_30_4966# VSUBS ground XM2/a_n50_n588# sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM3 ground ground ground ground VSUBS ground ground sky130_fd_pr__nfet_g5v0d10v5_NQCFE9
XXM4 ground ground ground ground VSUBS ground ground sky130_fd_pr__nfet_g5v0d10v5_CJGAEC
XXM5 m1_526_5878# m1_526_5878# m1_624_4748# m1_526_5878# m1_526_5878# m1_526_5878#
+ m1_526_5878# m1_526_5878# m1_526_5878# m1_624_4748# m1_624_4748# m1_624_4748# m1_624_4748#
+ m1_624_4748# m1_624_4748# m1_624_4748# m1_624_4748# m1_624_4748# m1_624_4748# m1_624_4748#
+ m1_624_4748# m1_624_4748# VSUBS m1_624_4748# m1_624_4748# sky130_fd_pr__nfet_g5v0d10v5_2MGL8M
XXM6 m1_n1264_7502# m1_n1222_6382# m1_n1264_7502# m1_n1264_7502# XM7/w_n586_n997#
+ m1_n1264_7502# m1_n1264_7502# m1_n1222_6382# m1_n1222_6382# m1_n1264_7502# sky130_fd_pr__pfet_g5v0d10v5_X3UTN5
XXM7 m1_62_6650# m1_n54_6380# m1_62_6650# m1_62_6650# XM7/w_n586_n997# m1_62_6650#
+ m1_62_6650# m1_n54_6380# m1_n54_6380# m1_62_6650# sky130_fd_pr__pfet_g5v0d10v5_AE43MT
XXM8 m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1458_8208#
+ m1_1458_8208# m1_1392_6382# m1_1392_6382# m1_1458_8208# m1_1458_8208# m1_1458_8208#
+ m1_1458_8208# m1_1392_6382# m1_1392_6382# m1_1392_6382# m1_1458_8208# m1_1458_8208#
+ m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1392_6382# m1_1392_6382# m1_1392_6382#
+ m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1392_6382#
+ m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1392_6382# m1_1392_6382# m1_1458_8208#
+ m1_1392_6382# m1_1392_6382# m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1392_6382#
+ m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1392_6382# m1_1458_8208# m1_1458_8208#
+ m1_1392_6382# m1_1392_6382# m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1392_6382#
+ m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1458_8208# m1_1392_6382# m1_1392_6382#
+ sky130_fd_pr__pfet_g5v0d10v5_CNRWF7
XXC1 sky130_fd_pr__cap_mim_m3_1_C5B489
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_C4MSH5 a_n69_630# a_n69_n1062# a_n199_n1192#
X0 a_n69_n1062# a_n69_630# a_n199_n1192# sky130_fd_pr__res_xhigh_po_0p69 l=6.3
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FG5HVM a_n100_n897# a_100_n800# a_n158_n800#
+ w_n358_n1097#
X0 a_100_n800# a_n100_n897# a_n158_n800# w_n358_n1097# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=2.32 ps=16.6 w=8 l=1
.ends

.subckt dac_cell4 vsup iref vsw iout iout_n vbias vgnd
XXR1 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69_C4MSH5
XXR2 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69_C4MSH5
XXR3 vsup parR vgnd sky130_fd_pr__res_xhigh_po_0p69_C4MSH5
XXR4 vsup parR vgnd sky130_fd_pr__res_xhigh_po_0p69_C4MSH5
XXM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5_FGUWVM
XXM2 iref sourceM3M4 sourceM2 vsup sky130_fd_pr__pfet_g5v0d10v5_FG5HVM
XXM3 vsw iout sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5_FG5HVM
XXM4 vbias iout_n sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5_FG5HVM
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_XZX24Q a_n199_n3262# a_n69_n3132# a_n69_2700#
X0 a_n69_n3132# a_n69_2700# a_n199_n3262# sky130_fd_pr__res_xhigh_po_0p69 l=27
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGK6VM a_n100_n297# a_100_n200# w_n358_n497#
+ a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n358_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt dac_cell2 vsup iref vsw iout iout_n vbias vgnd
XXR1 vgnd parR sourceM2 sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR2 vgnd parR sourceM2 sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR3 vgnd parR vsup sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR4 vgnd parR vsup sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5_FGUWVM
XXM2 iref sourceM3M4 vsup sourceM2 sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
XXM3 vsw iout vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
XXM4 vbias iout_n vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
.ends

.subckt dac_top_cell
Xdac_cell3_0 dac_cell3_0/vsup dac_cell3_0/iref dac_cell3_0/vsw dac_cell3_0/iout dac_cell3_0/iout_n
+ dac_cell3_0/vbias VSUBS dac_cell3
Xdac_cell1_0 dac_cell1_0/vsup dac_cell1_0/iref dac_cell1_0/vsw dac_cell1_0/iout dac_cell1_0/iout_n
+ dac_cell1_0/vbias VSUBS dac_cell1
Xmiel21_opamp_0 miel21_opamp_0/inPos miel21_opamp_0/inNeg miel21_opamp_0/outSingle
+ miel21_opamp_0/power miel21_opamp_0/ground VSUBS miel21_opamp
Xdac_cell4_0 dac_cell4_0/vsup dac_cell4_0/iref dac_cell4_0/vsw dac_cell4_0/iout dac_cell4_0/iout_n
+ dac_cell4_0/vbias VSUBS dac_cell4
Xdac_cell2_0 dac_cell2_0/vsup dac_cell2_0/iref dac_cell2_0/vsw dac_cell2_0/iout dac_cell2_0/iout_n
+ dac_cell2_0/vbias VSUBS dac_cell2
.ends

