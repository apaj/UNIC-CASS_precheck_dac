**.subckt opamp
V1 net1 GND 1
V2 net2 GND 1
V3 net3 GND 1
V4 net4 GND 1
XR1 net1 vin GND sky130_fd_pr__res_xhigh_po_5p73 L=2.8 mult=1 m=1
XR2 vin net2 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.8 mult=1 m=1
XR3 vin net3 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.8 mult=1 m=1
XR4 vin net4 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.8 mult=1 m=1
XR5 vin vout GND sky130_fd_pr__res_xhigh_po_5p73 L=2.8 mult=1 m=1
E1 vout GND vin GND 20000
**** begin user architecture code


.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.param mc_pr_switch=0
*** ANALYSIS TO DO

.tran 1m 100ms
.save 

.control
set wr_vecnames
set wr_singlescale


run
******** results filename  ************ nodes to write
***wrdata trans_opamp.res
.endc


**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.save
.end
