* SPICE3 file created from dac.ext - technology: sky130A

.subckt dac vdd vbias iout_neg iout vsw iin
X0 vdd vdd vdd sky130_fd_pr__res_iso_pw w=1.736e+07u l=1.325e+07u
X1 vdd vdd vdd sky130_fd_pr__res_iso_pw w=1.736e+07u l=1.325e+07u
X2 vdd vdd vdd sky130_fd_pr__res_iso_pw w=1.736e+07u l=1.325e+07u
X3 vdd vdd vdd sky130_fd_pr__res_iso_pw w=1.736e+07u l=1.325e+07u
X4 iin iin vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=1e+06u
X5 m1_1312_n646# iin vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6 iout_neg vbias m1_1312_n646# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X7 iout vsw m1_1312_n646# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
C0 vdd VSUBS 119.83fF
.ends
