magic
tech sky130A
timestamp 1698012353
use dac_top_cell  dac_top_cell_0 layout
timestamp 1698012353
transform 1 0 12271 0 1 9577
box -7190 -10182 12966 9172
<< end >>
