magic
tech sky130A
timestamp 1695294858
use top_dac  top_dac_0
timestamp 1695288709
transform 1 0 7068 0 1 -9
box 0 0 68000 84000
<< end >>
