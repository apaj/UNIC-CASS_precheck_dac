* SPICE3 file created from dac_cell3.ext - technology: sky130A

.option scale=5000u

.subckt dac_cell3 vsup vgnd iref vsw iout iout_n vbias
X0 m1_378_2344# li_n3490_2534# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=2600
X1 m1_378_2344# li_n3490_2534# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=2600
X2 vsup m1_378_2344# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=2600
X3 m1_378_2344# vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=2600
X4 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 ad=11600 pd=516 as=150800 ps=5664 w=200 l=200
X5 vsup iref li_n3490_2534# vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=800 l=200
X6 iout vsw vsup vsup sky130_fd_pr__pfet_g5v0d10v5 ad=46400 pd=1716 as=0 ps=0 w=800 l=200
X7 iout_n vbias vsup vsup sky130_fd_pr__pfet_g5v0d10v5 ad=46400 pd=1716 as=0 ps=0 w=800 l=200
.ends
