* NGSPICE file created from miel21_opamp.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p69_5CVACY a_n199_n1162# a_n69_600# a_n69_n1032#
X0 a_n69_600# a_n69_n1032# a_n199_n1162# sky130_fd_pr__res_xhigh_po_0p69 l=6
C0 a_n69_n1032# a_n199_n1162# 0.796f
C1 a_n69_600# a_n199_n1162# 0.796f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y a_50_n500# a_n242_n722# a_n108_n500# a_n50_n588#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n242_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
C0 a_n108_n500# a_50_n500# 0.562f
C1 a_50_n500# a_n242_n722# 0.61f
C2 a_n108_n500# a_n242_n722# 0.61f
C3 a_n50_n588# a_n242_n722# 0.455f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NQCFE9 a_189_n500# a_89_n588# a_31_n500# a_n189_n588#
+ a_n381_n722# a_n89_n500# a_n247_n500#
X0 a_189_n500# a_89_n588# a_31_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
X1 a_n89_n500# a_n189_n588# a_n247_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
C0 a_31_n500# a_189_n500# 0.562f
C1 a_31_n500# a_n89_n500# 0.833f
C2 a_n89_n500# a_n247_n500# 0.562f
C3 a_189_n500# a_n381_n722# 0.61f
C4 a_31_n500# a_n381_n722# 0.125f
C5 a_n89_n500# a_n381_n722# 0.125f
C6 a_n247_n500# a_n381_n722# 0.61f
C7 a_89_n588# a_n381_n722# 0.413f
C8 a_n189_n588# a_n381_n722# 0.413f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CJGAEC a_189_n500# a_89_n588# a_31_n500# a_n189_n588#
+ a_n381_n722# a_n89_n500# a_n247_n500#
X0 a_189_n500# a_89_n588# a_31_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
X1 a_n89_n500# a_n189_n588# a_n247_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
C0 a_31_n500# a_189_n500# 0.562f
C1 a_31_n500# a_n89_n500# 0.833f
C2 a_n89_n500# a_n247_n500# 0.562f
C3 a_189_n500# a_n381_n722# 0.61f
C4 a_31_n500# a_n381_n722# 0.125f
C5 a_n89_n500# a_n381_n722# 0.125f
C6 a_n247_n500# a_n381_n722# 0.61f
C7 a_89_n588# a_n381_n722# 0.413f
C8 a_n189_n588# a_n381_n722# 0.413f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2MGL8M a_367_n688# a_89_n688# a_31_n600# a_n189_n688#
+ a_n1023_n688# a_645_n688# a_n467_n688# a_923_n688# a_n745_n688# a_n89_n600# a_n367_n600#
+ a_n645_n600# a_n1081_n600# a_n247_n600# a_n923_n600# a_n525_n600# a_n803_n600# a_309_n600#
+ a_587_n600# a_189_n600# a_865_n600# a_467_n600# a_n1215_n822# a_745_n600# a_1023_n600#
X0 a_n367_n600# a_n467_n688# a_n525_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X1 a_467_n600# a_367_n688# a_309_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X2 a_189_n600# a_89_n688# a_31_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X3 a_n645_n600# a_n745_n688# a_n803_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X4 a_745_n600# a_645_n688# a_587_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X5 a_n89_n600# a_n189_n688# a_n247_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X6 a_n923_n600# a_n1023_n688# a_n1081_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X7 a_1023_n600# a_923_n688# a_865_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
C0 a_745_n600# a_865_n600# 0.999f
C1 a_n923_n600# a_n803_n600# 0.999f
C2 a_n367_n600# a_n247_n600# 0.999f
C3 a_n89_n600# a_31_n600# 0.999f
C4 a_467_n600# a_587_n600# 0.999f
C5 a_1023_n600# a_865_n600# 0.674f
C6 a_n89_n600# a_n247_n600# 0.674f
C7 a_189_n600# a_309_n600# 0.999f
C8 a_n525_n600# a_n367_n600# 0.674f
C9 a_n803_n600# a_n645_n600# 0.674f
C10 a_745_n600# a_587_n600# 0.674f
C11 a_309_n600# a_467_n600# 0.674f
C12 a_n923_n600# a_n1081_n600# 0.674f
C13 a_189_n600# a_31_n600# 0.674f
C14 a_n525_n600# a_n645_n600# 0.999f
C15 a_1023_n600# a_n1215_n822# 0.725f
C16 a_865_n600# a_n1215_n822# 0.143f
C17 a_745_n600# a_n1215_n822# 0.143f
C18 a_587_n600# a_n1215_n822# 0.143f
C19 a_467_n600# a_n1215_n822# 0.143f
C20 a_309_n600# a_n1215_n822# 0.143f
C21 a_189_n600# a_n1215_n822# 0.143f
C22 a_31_n600# a_n1215_n822# 0.143f
C23 a_n89_n600# a_n1215_n822# 0.143f
C24 a_n247_n600# a_n1215_n822# 0.143f
C25 a_n367_n600# a_n1215_n822# 0.143f
C26 a_n525_n600# a_n1215_n822# 0.143f
C27 a_n645_n600# a_n1215_n822# 0.143f
C28 a_n803_n600# a_n1215_n822# 0.143f
C29 a_n923_n600# a_n1215_n822# 0.143f
C30 a_n1081_n600# a_n1215_n822# 0.725f
C31 a_923_n688# a_n1215_n822# 0.414f
C32 a_645_n688# a_n1215_n822# 0.371f
C33 a_367_n688# a_n1215_n822# 0.371f
C34 a_89_n688# a_n1215_n822# 0.371f
C35 a_n189_n688# a_n1215_n822# 0.371f
C36 a_n467_n688# a_n1215_n822# 0.371f
C37 a_n745_n688# a_n1215_n822# 0.371f
C38 a_n1023_n688# a_n1215_n822# 0.414f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_X3UTN5 a_170_n700# a_n50_n797# a_50_n700# a_n228_n700#
+ w_n586_n997# a_n108_n700# a_n386_n700# a_228_n797# a_n328_n797# a_328_n700# VSUBS
X0 a_328_n700# a_228_n797# a_170_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X1 a_50_n700# a_n50_n797# a_n108_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X2 a_n228_n700# a_n328_n797# a_n386_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
C0 a_228_n797# w_n586_n997# 0.111f
C1 w_n586_n997# a_328_n700# 0.534f
C2 a_n228_n700# a_n386_n700# 0.786f
C3 w_n586_n997# a_n386_n700# 0.534f
C4 a_170_n700# a_328_n700# 0.786f
C5 a_170_n700# a_50_n700# 1.16f
C6 w_n586_n997# a_n328_n797# 0.111f
C7 a_n108_n700# a_50_n700# 0.786f
C8 a_n228_n700# a_n108_n700# 1.16f
C9 a_328_n700# VSUBS 0.308f
C10 a_170_n700# VSUBS 0.106f
C11 a_50_n700# VSUBS 0.106f
C12 a_n108_n700# VSUBS 0.106f
C13 a_n228_n700# VSUBS 0.106f
C14 a_n386_n700# VSUBS 0.308f
C15 a_228_n797# VSUBS 0.148f
C16 a_n50_n797# VSUBS 0.124f
C17 a_n328_n797# VSUBS 0.148f
C18 w_n586_n997# VSUBS 8.51f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AE43MT a_170_n700# a_n50_n797# a_50_n700# a_n228_n700#
+ w_n586_n997# a_n108_n700# a_n386_n700# a_228_n797# a_n328_n797# a_328_n700# VSUBS
X0 a_328_n700# a_228_n797# a_170_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X1 a_50_n700# a_n50_n797# a_n108_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X2 a_n228_n700# a_n328_n797# a_n386_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
C0 a_50_n700# a_n108_n700# 0.786f
C1 w_n586_n997# a_n386_n700# 0.534f
C2 w_n586_n997# a_328_n700# 0.534f
C3 a_n386_n700# a_n228_n700# 0.786f
C4 w_n586_n997# a_228_n797# 0.111f
C5 a_n108_n700# a_n228_n700# 1.16f
C6 w_n586_n997# a_n328_n797# 0.111f
C7 a_50_n700# a_170_n700# 1.16f
C8 a_170_n700# a_328_n700# 0.786f
C9 a_328_n700# VSUBS 0.308f
C10 a_170_n700# VSUBS 0.106f
C11 a_50_n700# VSUBS 0.106f
C12 a_n108_n700# VSUBS 0.106f
C13 a_n228_n700# VSUBS 0.106f
C14 a_n386_n700# VSUBS 0.308f
C15 a_228_n797# VSUBS 0.148f
C16 a_n50_n797# VSUBS 0.124f
C17 a_n328_n797# VSUBS 0.148f
C18 w_n586_n997# VSUBS 8.51f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CNRWF7 a_1579_n1300# a_n803_n1300# a_n1757_n1300#
+ a_n2035_n1300# a_1301_n1300# a_n645_n1300# a_1143_n1300# a_n2413_n1397# a_n2691_n1397#
+ a_n1637_n1300# a_n2193_n1300# w_n2949_n1597# a_189_n1300# a_n525_n1300# a_2591_n1397#
+ a_2313_n1397# a_923_n1397# a_2533_n1300# a_1023_n1300# a_n1479_n1300# a_n367_n1300#
+ a_n1201_n1300# a_n1857_n1397# a_n2135_n1397# a_n745_n1397# a_2691_n1300# a_2413_n1300#
+ a_n89_n1300# a_n1359_n1300# a_n247_n1300# a_645_n1397# a_2255_n1300# a_1977_n1300#
+ a_865_n1300# a_2035_n1397# a_1757_n1397# a_n2749_n1300# a_n1579_n1397# a_n1301_n1397#
+ a_2135_n1300# a_1857_n1300# a_745_n1300# a_n467_n1397# a_n1081_n1300# a_n2313_n1300#
+ a_n2591_n1300# a_89_n1397# a_587_n1300# a_309_n1300# a_1479_n1397# a_367_n1397#
+ a_1699_n1300# a_31_n1300# a_n923_n1300# a_1201_n1397# a_1421_n1300# a_n1915_n1300#
+ a_n2471_n1300# a_467_n1300# a_n189_n1397# a_n1023_n1397# VSUBS
X0 a_1857_n1300# a_1757_n1397# a_1699_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X1 a_2691_n1300# a_2591_n1397# a_2533_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X2 a_n923_n1300# a_n1023_n1397# a_n1081_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X3 a_745_n1300# a_645_n1397# a_587_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X4 a_n2035_n1300# a_n2135_n1397# a_n2193_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X5 a_1579_n1300# a_1479_n1397# a_1421_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X6 a_467_n1300# a_367_n1397# a_309_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X7 a_n645_n1300# a_n745_n1397# a_n803_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X8 a_n2591_n1300# a_n2691_n1397# a_n2749_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X9 a_n1757_n1300# a_n1857_n1397# a_n1915_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X10 a_n367_n1300# a_n467_n1397# a_n525_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X11 a_1301_n1300# a_1201_n1397# a_1143_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X12 a_2413_n1300# a_2313_n1397# a_2255_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X13 a_n1479_n1300# a_n1579_n1397# a_n1637_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X14 a_n89_n1300# a_n189_n1397# a_n247_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X15 a_2135_n1300# a_2035_n1397# a_1977_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X16 a_189_n1300# a_89_n1397# a_31_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X17 a_n1201_n1300# a_n1301_n1397# a_n1359_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X18 a_1023_n1300# a_923_n1397# a_865_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X19 a_n2313_n1300# a_n2413_n1397# a_n2471_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
C0 a_n2691_n1397# w_n2949_n1597# 0.111f
C1 a_n923_n1300# a_n1023_n1397# 0.165f
C2 a_865_n1300# a_745_n1300# 2.16f
C3 a_189_n1300# a_309_n1300# 2.16f
C4 a_865_n1300# a_1023_n1300# 1.46f
C5 a_n745_n1397# a_n803_n1300# 0.165f
C6 a_n189_n1397# a_n89_n1300# 0.165f
C7 a_n923_n1300# a_n1081_n1300# 1.46f
C8 a_2413_n1300# a_2313_n1397# 0.165f
C9 a_n1359_n1300# a_n1479_n1300# 2.16f
C10 a_n2691_n1397# a_n2749_n1300# 0.165f
C11 a_1857_n1300# a_1977_n1300# 2.16f
C12 a_1757_n1397# a_1857_n1300# 0.165f
C13 a_2255_n1300# a_2413_n1300# 1.46f
C14 a_n2035_n1300# a_n2135_n1397# 0.165f
C15 a_n247_n1300# a_n367_n1300# 2.16f
C16 a_n1757_n1300# a_n1637_n1300# 2.16f
C17 a_1757_n1397# a_1699_n1300# 0.165f
C18 a_n2749_n1300# a_n2591_n1300# 1.46f
C19 a_n247_n1300# a_n89_n1300# 1.46f
C20 a_1421_n1300# a_1579_n1300# 1.46f
C21 a_2255_n1300# a_2313_n1397# 0.165f
C22 a_2035_n1397# a_2135_n1300# 0.165f
C23 a_n1637_n1300# a_n1479_n1300# 1.46f
C24 a_n1201_n1300# a_n1081_n1300# 2.16f
C25 a_2413_n1300# a_2533_n1300# 2.16f
C26 a_1023_n1300# a_1143_n1300# 2.16f
C27 a_1977_n1300# a_2035_n1397# 0.165f
C28 a_n525_n1300# a_n367_n1300# 1.46f
C29 a_n2413_n1397# a_n2471_n1300# 0.165f
C30 a_n923_n1300# a_n803_n1300# 2.16f
C31 a_n1081_n1300# a_n1023_n1397# 0.165f
C32 a_1201_n1397# a_1143_n1300# 0.165f
C33 a_645_n1397# a_587_n1300# 0.165f
C34 a_n1757_n1300# a_n1915_n1300# 1.46f
C35 a_n525_n1300# a_n645_n1300# 2.16f
C36 a_n645_n1300# a_n803_n1300# 1.46f
C37 a_n2471_n1300# a_n2313_n1300# 1.46f
C38 a_n2591_n1300# a_n2471_n1300# 2.16f
C39 a_n1757_n1300# a_n1857_n1397# 0.165f
C40 a_n525_n1300# a_n467_n1397# 0.165f
C41 a_367_n1397# a_467_n1300# 0.165f
C42 a_n2749_n1300# w_n2949_n1597# 0.967f
C43 a_n1359_n1300# a_n1201_n1300# 1.46f
C44 a_n2035_n1300# a_n1915_n1300# 2.16f
C45 a_n745_n1397# a_n645_n1300# 0.165f
C46 a_n1201_n1300# a_n1301_n1397# 0.165f
C47 a_1977_n1300# a_2135_n1300# 1.46f
C48 a_n247_n1300# a_n189_n1397# 0.165f
C49 a_31_n1300# a_89_n1397# 0.165f
C50 a_1421_n1300# a_1479_n1397# 0.165f
C51 w_n2949_n1597# a_2591_n1397# 0.111f
C52 a_467_n1300# a_587_n1300# 2.16f
C53 a_367_n1397# a_309_n1300# 0.165f
C54 a_n2413_n1397# a_n2313_n1300# 0.165f
C55 a_n2193_n1300# a_n2313_n1300# 2.16f
C56 a_2691_n1300# w_n2949_n1597# 0.967f
C57 a_865_n1300# a_923_n1397# 0.165f
C58 a_1201_n1397# a_1301_n1300# 0.165f
C59 a_n2691_n1397# a_n2591_n1300# 0.165f
C60 a_1579_n1300# a_1699_n1300# 2.16f
C61 a_1857_n1300# a_1699_n1300# 1.46f
C62 a_2533_n1300# a_2591_n1397# 0.165f
C63 a_n89_n1300# a_31_n1300# 2.16f
C64 a_189_n1300# a_89_n1397# 0.165f
C65 a_n1857_n1397# a_n1915_n1300# 0.165f
C66 a_645_n1397# a_745_n1300# 0.165f
C67 a_1143_n1300# a_1301_n1300# 1.46f
C68 a_n2193_n1300# a_n2135_n1397# 0.165f
C69 a_923_n1397# a_1023_n1300# 0.165f
C70 a_587_n1300# a_745_n1300# 1.46f
C71 a_n367_n1300# a_n467_n1397# 0.165f
C72 a_2691_n1300# a_2533_n1300# 1.46f
C73 a_189_n1300# a_31_n1300# 1.46f
C74 a_n1579_n1397# a_n1637_n1300# 0.165f
C75 a_2255_n1300# a_2135_n1300# 2.16f
C76 a_309_n1300# a_467_n1300# 1.46f
C77 a_n1359_n1300# a_n1301_n1397# 0.165f
C78 a_2691_n1300# a_2591_n1397# 0.165f
C79 a_n1579_n1397# a_n1479_n1300# 0.165f
C80 a_n2193_n1300# a_n2035_n1300# 1.46f
C81 a_1479_n1397# a_1579_n1300# 0.165f
C82 a_1421_n1300# a_1301_n1300# 2.16f
C83 a_2691_n1300# VSUBS 0.565f
C84 a_2533_n1300# VSUBS 0.19f
C85 a_2413_n1300# VSUBS 0.19f
C86 a_2255_n1300# VSUBS 0.19f
C87 a_2135_n1300# VSUBS 0.19f
C88 a_1977_n1300# VSUBS 0.19f
C89 a_1857_n1300# VSUBS 0.19f
C90 a_1699_n1300# VSUBS 0.19f
C91 a_1579_n1300# VSUBS 0.19f
C92 a_1421_n1300# VSUBS 0.19f
C93 a_1301_n1300# VSUBS 0.19f
C94 a_1143_n1300# VSUBS 0.19f
C95 a_1023_n1300# VSUBS 0.19f
C96 a_865_n1300# VSUBS 0.19f
C97 a_745_n1300# VSUBS 0.19f
C98 a_587_n1300# VSUBS 0.19f
C99 a_467_n1300# VSUBS 0.19f
C100 a_309_n1300# VSUBS 0.19f
C101 a_189_n1300# VSUBS 0.19f
C102 a_31_n1300# VSUBS 0.19f
C103 a_n89_n1300# VSUBS 0.19f
C104 a_n247_n1300# VSUBS 0.19f
C105 a_n367_n1300# VSUBS 0.19f
C106 a_n525_n1300# VSUBS 0.19f
C107 a_n645_n1300# VSUBS 0.19f
C108 a_n803_n1300# VSUBS 0.19f
C109 a_n923_n1300# VSUBS 0.19f
C110 a_n1081_n1300# VSUBS 0.19f
C111 a_n1201_n1300# VSUBS 0.19f
C112 a_n1359_n1300# VSUBS 0.19f
C113 a_n1479_n1300# VSUBS 0.19f
C114 a_n1637_n1300# VSUBS 0.19f
C115 a_n1757_n1300# VSUBS 0.19f
C116 a_n1915_n1300# VSUBS 0.19f
C117 a_n2035_n1300# VSUBS 0.19f
C118 a_n2193_n1300# VSUBS 0.19f
C119 a_n2313_n1300# VSUBS 0.19f
C120 a_n2471_n1300# VSUBS 0.19f
C121 a_n2591_n1300# VSUBS 0.19f
C122 a_n2749_n1300# VSUBS 0.565f
C123 a_2591_n1397# VSUBS 0.159f
C124 a_2313_n1397# VSUBS 0.136f
C125 a_2035_n1397# VSUBS 0.136f
C126 a_1757_n1397# VSUBS 0.136f
C127 a_1479_n1397# VSUBS 0.136f
C128 a_1201_n1397# VSUBS 0.136f
C129 a_923_n1397# VSUBS 0.136f
C130 a_645_n1397# VSUBS 0.136f
C131 a_367_n1397# VSUBS 0.136f
C132 a_89_n1397# VSUBS 0.136f
C133 a_n189_n1397# VSUBS 0.136f
C134 a_n467_n1397# VSUBS 0.136f
C135 a_n745_n1397# VSUBS 0.136f
C136 a_n1023_n1397# VSUBS 0.136f
C137 a_n1301_n1397# VSUBS 0.136f
C138 a_n1579_n1397# VSUBS 0.136f
C139 a_n1857_n1397# VSUBS 0.136f
C140 a_n2135_n1397# VSUBS 0.136f
C141 a_n2413_n1397# VSUBS 0.136f
C142 a_n2691_n1397# VSUBS 0.159f
C143 w_n2949_n1597# VSUBS 61.7f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_C5B489 c1_n1050_n1400# m3_n1150_n1500# VSUBS
X0 c1_n1050_n1400# m3_n1150_n1500# sky130_fd_pr__cap_mim_m3_1 l=14 w=10
C0 m3_n1150_n1500# c1_n1050_n1400# 14f
C1 c1_n1050_n1400# VSUBS 1.11f
C2 m3_n1150_n1500# VSUBS 4.9f
.ends

.subckt miel21_opamp inPos inNeg outSingle power ground
XXR1 ground m1_n1838_8400# bias sky130_fd_pr__res_xhigh_po_0p69_5CVACY
XXR2 ground m1_n1838_8400# m1_360_8394# sky130_fd_pr__res_xhigh_po_0p69_5CVACY
XXR3 ground m1_360_8394# power sky130_fd_pr__res_xhigh_po_0p69_5CVACY
XXM1 d1 ground nsources inPos sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM2 d2 ground nsources inNeg sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM3 bias bias ground bias ground bias ground sky130_fd_pr__nfet_g5v0d10v5_NQCFE9
XXM4 nsources bias ground bias ground nsources ground sky130_fd_pr__nfet_g5v0d10v5_CJGAEC
XXM5 bias bias ground bias bias bias bias bias bias outSingle outSingle outSingle
+ ground ground outSingle ground ground ground ground outSingle ground outSingle ground
+ outSingle outSingle sky130_fd_pr__nfet_g5v0d10v5_2MGL8M
XXM6 power d1 d1 d1 power power power d1 d1 d1 ground sky130_fd_pr__pfet_g5v0d10v5_X3UTN5
XXM7 power d1 d2 d2 power power power d1 d1 d2 ground sky130_fd_pr__pfet_g5v0d10v5_AE43MT
XXM8 outSingle power outSingle outSingle outSingle outSingle power d2 d2 power power
+ power outSingle power d2 d2 d2 power outSingle outSingle outSingle outSingle d2
+ d2 d2 outSingle outSingle outSingle power power d2 power power power d2 d2 power
+ d2 d2 outSingle outSingle outSingle d2 power outSingle outSingle d2 power power
+ d2 d2 power power outSingle d2 power power power outSingle d2 d2 ground sky130_fd_pr__pfet_g5v0d10v5_CNRWF7
XXC1 outSingle d2 ground sky130_fd_pr__cap_mim_m3_1_C5B489
C0 m1_n1838_8400# power 0.268f
C1 inPos bias 0.532f
C2 bias d2 0.146f
C3 m1_360_8394# power 0.249f
C4 nsources d1 1.13f
C5 bias power 0.19f
C6 d2 power 7.01f
C7 inNeg nsources 0.268f
C8 outSingle bias 1.15f
C9 outSingle d2 4.44f
C10 outSingle power 10.3f
C11 bias d1 0.368f
C12 inPos d1 0.12f
C13 d1 d2 0.545f
C14 bias nsources 0.394f
C15 inPos nsources 0.129f
C16 nsources d2 0.201f
C17 nsources m1_n126_4512# 0.109f
C18 d1 power 3.18f
C19 inNeg bias 1.06f
C20 inNeg inPos 0.596f
C21 m1_n126_4512# ground 0.135f $ **FLOATING
C22 power ground 85.9f
C23 outSingle ground 14.8f
C24 nsources ground 3.29f
C25 bias ground 15.2f
C26 d2 ground 11.1f
C27 inNeg ground 1.98f
C28 d1 ground 2.32f
C29 inPos ground 2.85f
C30 m1_360_8394# ground 1.64f
C31 m1_n1838_8400# ground 2.1f
.ends

