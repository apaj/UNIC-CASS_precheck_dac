magic
tech sky130A
magscale 1 2
timestamp 1697533315
<< pwell >>
rect -357 -758 357 758
<< mvnmos >>
rect -129 -500 -29 500
rect 29 -500 129 500
<< mvndiff >>
rect -187 488 -129 500
rect -187 -488 -175 488
rect -141 -488 -129 488
rect -187 -500 -129 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 129 488 187 500
rect 129 -488 141 488
rect 175 -488 187 488
rect 129 -500 187 -488
<< mvndiffc >>
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
<< mvpsubdiff >>
rect -321 710 321 722
rect -321 676 -213 710
rect 213 676 321 710
rect -321 664 321 676
rect -321 614 -263 664
rect -321 -614 -309 614
rect -275 -614 -263 614
rect 263 614 321 664
rect -321 -664 -263 -614
rect 263 -614 275 614
rect 309 -614 321 614
rect 263 -664 321 -614
rect -321 -676 321 -664
rect -321 -710 -213 -676
rect 213 -710 321 -676
rect -321 -722 321 -710
<< mvpsubdiffcont >>
rect -213 676 213 710
rect -309 -614 -275 614
rect 275 -614 309 614
rect -213 -710 213 -676
<< poly >>
rect -129 572 -29 588
rect -129 538 -113 572
rect -45 538 -29 572
rect -129 500 -29 538
rect 29 572 129 588
rect 29 538 45 572
rect 113 538 129 572
rect 29 500 129 538
rect -129 -538 -29 -500
rect -129 -572 -113 -538
rect -45 -572 -29 -538
rect -129 -588 -29 -572
rect 29 -538 129 -500
rect 29 -572 45 -538
rect 113 -572 129 -538
rect 29 -588 129 -572
<< polycont >>
rect -113 538 -45 572
rect 45 538 113 572
rect -113 -572 -45 -538
rect 45 -572 113 -538
<< locali >>
rect -309 676 -213 710
rect 213 676 309 710
rect -309 614 -275 676
rect 275 614 309 676
rect -129 538 -113 572
rect -45 538 -29 572
rect 29 538 45 572
rect 113 538 129 572
rect -175 488 -141 504
rect -175 -504 -141 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 141 488 175 504
rect 141 -504 175 -488
rect -129 -572 -113 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 113 -572 129 -538
rect -309 -676 -275 -614
rect 275 -676 309 -614
rect -309 -710 -213 -676
rect 213 -710 309 -676
<< viali >>
rect -113 538 -45 572
rect 45 538 113 572
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect -113 -572 -45 -538
rect 45 -572 113 -538
<< metal1 >>
rect -125 572 -33 578
rect -125 538 -113 572
rect -45 538 -33 572
rect -125 532 -33 538
rect 33 572 125 578
rect 33 538 45 572
rect 113 538 125 572
rect 33 532 125 538
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -181 -500 -135 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 135 488 181 500
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect -125 -538 -33 -532
rect -125 -572 -113 -538
rect -45 -572 -33 -538
rect -125 -578 -33 -572
rect 33 -538 125 -532
rect 33 -572 45 -538
rect 113 -572 125 -538
rect 33 -578 125 -572
<< properties >>
string FIXED_BBOX -292 -693 292 693
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
