magic
tech sky130A
magscale 1 2
timestamp 1696876712
<< nwell >>
rect -925 -1269 925 1269
<< mvpmos >>
rect -667 772 -467 972
rect -289 772 -89 972
rect 89 772 289 972
rect 467 772 667 972
rect -667 336 -467 536
rect -289 336 -89 536
rect 89 336 289 536
rect 467 336 667 536
rect -667 -100 -467 100
rect -289 -100 -89 100
rect 89 -100 289 100
rect 467 -100 667 100
rect -667 -536 -467 -336
rect -289 -536 -89 -336
rect 89 -536 289 -336
rect 467 -536 667 -336
rect -667 -972 -467 -772
rect -289 -972 -89 -772
rect 89 -972 289 -772
rect 467 -972 667 -772
<< mvpdiff >>
rect -725 960 -667 972
rect -725 784 -713 960
rect -679 784 -667 960
rect -725 772 -667 784
rect -467 960 -409 972
rect -467 784 -455 960
rect -421 784 -409 960
rect -467 772 -409 784
rect -347 960 -289 972
rect -347 784 -335 960
rect -301 784 -289 960
rect -347 772 -289 784
rect -89 960 -31 972
rect -89 784 -77 960
rect -43 784 -31 960
rect -89 772 -31 784
rect 31 960 89 972
rect 31 784 43 960
rect 77 784 89 960
rect 31 772 89 784
rect 289 960 347 972
rect 289 784 301 960
rect 335 784 347 960
rect 289 772 347 784
rect 409 960 467 972
rect 409 784 421 960
rect 455 784 467 960
rect 409 772 467 784
rect 667 960 725 972
rect 667 784 679 960
rect 713 784 725 960
rect 667 772 725 784
rect -725 524 -667 536
rect -725 348 -713 524
rect -679 348 -667 524
rect -725 336 -667 348
rect -467 524 -409 536
rect -467 348 -455 524
rect -421 348 -409 524
rect -467 336 -409 348
rect -347 524 -289 536
rect -347 348 -335 524
rect -301 348 -289 524
rect -347 336 -289 348
rect -89 524 -31 536
rect -89 348 -77 524
rect -43 348 -31 524
rect -89 336 -31 348
rect 31 524 89 536
rect 31 348 43 524
rect 77 348 89 524
rect 31 336 89 348
rect 289 524 347 536
rect 289 348 301 524
rect 335 348 347 524
rect 289 336 347 348
rect 409 524 467 536
rect 409 348 421 524
rect 455 348 467 524
rect 409 336 467 348
rect 667 524 725 536
rect 667 348 679 524
rect 713 348 725 524
rect 667 336 725 348
rect -725 88 -667 100
rect -725 -88 -713 88
rect -679 -88 -667 88
rect -725 -100 -667 -88
rect -467 88 -409 100
rect -467 -88 -455 88
rect -421 -88 -409 88
rect -467 -100 -409 -88
rect -347 88 -289 100
rect -347 -88 -335 88
rect -301 -88 -289 88
rect -347 -100 -289 -88
rect -89 88 -31 100
rect -89 -88 -77 88
rect -43 -88 -31 88
rect -89 -100 -31 -88
rect 31 88 89 100
rect 31 -88 43 88
rect 77 -88 89 88
rect 31 -100 89 -88
rect 289 88 347 100
rect 289 -88 301 88
rect 335 -88 347 88
rect 289 -100 347 -88
rect 409 88 467 100
rect 409 -88 421 88
rect 455 -88 467 88
rect 409 -100 467 -88
rect 667 88 725 100
rect 667 -88 679 88
rect 713 -88 725 88
rect 667 -100 725 -88
rect -725 -348 -667 -336
rect -725 -524 -713 -348
rect -679 -524 -667 -348
rect -725 -536 -667 -524
rect -467 -348 -409 -336
rect -467 -524 -455 -348
rect -421 -524 -409 -348
rect -467 -536 -409 -524
rect -347 -348 -289 -336
rect -347 -524 -335 -348
rect -301 -524 -289 -348
rect -347 -536 -289 -524
rect -89 -348 -31 -336
rect -89 -524 -77 -348
rect -43 -524 -31 -348
rect -89 -536 -31 -524
rect 31 -348 89 -336
rect 31 -524 43 -348
rect 77 -524 89 -348
rect 31 -536 89 -524
rect 289 -348 347 -336
rect 289 -524 301 -348
rect 335 -524 347 -348
rect 289 -536 347 -524
rect 409 -348 467 -336
rect 409 -524 421 -348
rect 455 -524 467 -348
rect 409 -536 467 -524
rect 667 -348 725 -336
rect 667 -524 679 -348
rect 713 -524 725 -348
rect 667 -536 725 -524
rect -725 -784 -667 -772
rect -725 -960 -713 -784
rect -679 -960 -667 -784
rect -725 -972 -667 -960
rect -467 -784 -409 -772
rect -467 -960 -455 -784
rect -421 -960 -409 -784
rect -467 -972 -409 -960
rect -347 -784 -289 -772
rect -347 -960 -335 -784
rect -301 -960 -289 -784
rect -347 -972 -289 -960
rect -89 -784 -31 -772
rect -89 -960 -77 -784
rect -43 -960 -31 -784
rect -89 -972 -31 -960
rect 31 -784 89 -772
rect 31 -960 43 -784
rect 77 -960 89 -784
rect 31 -972 89 -960
rect 289 -784 347 -772
rect 289 -960 301 -784
rect 335 -960 347 -784
rect 289 -972 347 -960
rect 409 -784 467 -772
rect 409 -960 421 -784
rect 455 -960 467 -784
rect 409 -972 467 -960
rect 667 -784 725 -772
rect 667 -960 679 -784
rect 713 -960 725 -784
rect 667 -972 725 -960
<< mvpdiffc >>
rect -713 784 -679 960
rect -455 784 -421 960
rect -335 784 -301 960
rect -77 784 -43 960
rect 43 784 77 960
rect 301 784 335 960
rect 421 784 455 960
rect 679 784 713 960
rect -713 348 -679 524
rect -455 348 -421 524
rect -335 348 -301 524
rect -77 348 -43 524
rect 43 348 77 524
rect 301 348 335 524
rect 421 348 455 524
rect 679 348 713 524
rect -713 -88 -679 88
rect -455 -88 -421 88
rect -335 -88 -301 88
rect -77 -88 -43 88
rect 43 -88 77 88
rect 301 -88 335 88
rect 421 -88 455 88
rect 679 -88 713 88
rect -713 -524 -679 -348
rect -455 -524 -421 -348
rect -335 -524 -301 -348
rect -77 -524 -43 -348
rect 43 -524 77 -348
rect 301 -524 335 -348
rect 421 -524 455 -348
rect 679 -524 713 -348
rect -713 -960 -679 -784
rect -455 -960 -421 -784
rect -335 -960 -301 -784
rect -77 -960 -43 -784
rect 43 -960 77 -784
rect 301 -960 335 -784
rect 421 -960 455 -784
rect 679 -960 713 -784
<< mvnsubdiff >>
rect -859 1191 859 1203
rect -859 1157 -751 1191
rect 751 1157 859 1191
rect -859 1145 859 1157
rect -859 1095 -801 1145
rect -859 -1095 -847 1095
rect -813 -1095 -801 1095
rect 801 1095 859 1145
rect -859 -1145 -801 -1095
rect 801 -1095 813 1095
rect 847 -1095 859 1095
rect 801 -1145 859 -1095
rect -859 -1157 859 -1145
rect -859 -1191 -751 -1157
rect 751 -1191 859 -1157
rect -859 -1203 859 -1191
<< mvnsubdiffcont >>
rect -751 1157 751 1191
rect -847 -1095 -813 1095
rect 813 -1095 847 1095
rect -751 -1191 751 -1157
<< poly >>
rect -667 1053 -467 1069
rect -667 1019 -651 1053
rect -483 1019 -467 1053
rect -667 972 -467 1019
rect -289 1053 -89 1069
rect -289 1019 -273 1053
rect -105 1019 -89 1053
rect -289 972 -89 1019
rect 89 1053 289 1069
rect 89 1019 105 1053
rect 273 1019 289 1053
rect 89 972 289 1019
rect 467 1053 667 1069
rect 467 1019 483 1053
rect 651 1019 667 1053
rect 467 972 667 1019
rect -667 725 -467 772
rect -667 691 -651 725
rect -483 691 -467 725
rect -667 675 -467 691
rect -289 725 -89 772
rect -289 691 -273 725
rect -105 691 -89 725
rect -289 675 -89 691
rect 89 725 289 772
rect 89 691 105 725
rect 273 691 289 725
rect 89 675 289 691
rect 467 725 667 772
rect 467 691 483 725
rect 651 691 667 725
rect 467 675 667 691
rect -667 617 -467 633
rect -667 583 -651 617
rect -483 583 -467 617
rect -667 536 -467 583
rect -289 617 -89 633
rect -289 583 -273 617
rect -105 583 -89 617
rect -289 536 -89 583
rect 89 617 289 633
rect 89 583 105 617
rect 273 583 289 617
rect 89 536 289 583
rect 467 617 667 633
rect 467 583 483 617
rect 651 583 667 617
rect 467 536 667 583
rect -667 289 -467 336
rect -667 255 -651 289
rect -483 255 -467 289
rect -667 239 -467 255
rect -289 289 -89 336
rect -289 255 -273 289
rect -105 255 -89 289
rect -289 239 -89 255
rect 89 289 289 336
rect 89 255 105 289
rect 273 255 289 289
rect 89 239 289 255
rect 467 289 667 336
rect 467 255 483 289
rect 651 255 667 289
rect 467 239 667 255
rect -667 181 -467 197
rect -667 147 -651 181
rect -483 147 -467 181
rect -667 100 -467 147
rect -289 181 -89 197
rect -289 147 -273 181
rect -105 147 -89 181
rect -289 100 -89 147
rect 89 181 289 197
rect 89 147 105 181
rect 273 147 289 181
rect 89 100 289 147
rect 467 181 667 197
rect 467 147 483 181
rect 651 147 667 181
rect 467 100 667 147
rect -667 -147 -467 -100
rect -667 -181 -651 -147
rect -483 -181 -467 -147
rect -667 -197 -467 -181
rect -289 -147 -89 -100
rect -289 -181 -273 -147
rect -105 -181 -89 -147
rect -289 -197 -89 -181
rect 89 -147 289 -100
rect 89 -181 105 -147
rect 273 -181 289 -147
rect 89 -197 289 -181
rect 467 -147 667 -100
rect 467 -181 483 -147
rect 651 -181 667 -147
rect 467 -197 667 -181
rect -667 -255 -467 -239
rect -667 -289 -651 -255
rect -483 -289 -467 -255
rect -667 -336 -467 -289
rect -289 -255 -89 -239
rect -289 -289 -273 -255
rect -105 -289 -89 -255
rect -289 -336 -89 -289
rect 89 -255 289 -239
rect 89 -289 105 -255
rect 273 -289 289 -255
rect 89 -336 289 -289
rect 467 -255 667 -239
rect 467 -289 483 -255
rect 651 -289 667 -255
rect 467 -336 667 -289
rect -667 -583 -467 -536
rect -667 -617 -651 -583
rect -483 -617 -467 -583
rect -667 -633 -467 -617
rect -289 -583 -89 -536
rect -289 -617 -273 -583
rect -105 -617 -89 -583
rect -289 -633 -89 -617
rect 89 -583 289 -536
rect 89 -617 105 -583
rect 273 -617 289 -583
rect 89 -633 289 -617
rect 467 -583 667 -536
rect 467 -617 483 -583
rect 651 -617 667 -583
rect 467 -633 667 -617
rect -667 -691 -467 -675
rect -667 -725 -651 -691
rect -483 -725 -467 -691
rect -667 -772 -467 -725
rect -289 -691 -89 -675
rect -289 -725 -273 -691
rect -105 -725 -89 -691
rect -289 -772 -89 -725
rect 89 -691 289 -675
rect 89 -725 105 -691
rect 273 -725 289 -691
rect 89 -772 289 -725
rect 467 -691 667 -675
rect 467 -725 483 -691
rect 651 -725 667 -691
rect 467 -772 667 -725
rect -667 -1019 -467 -972
rect -667 -1053 -651 -1019
rect -483 -1053 -467 -1019
rect -667 -1069 -467 -1053
rect -289 -1019 -89 -972
rect -289 -1053 -273 -1019
rect -105 -1053 -89 -1019
rect -289 -1069 -89 -1053
rect 89 -1019 289 -972
rect 89 -1053 105 -1019
rect 273 -1053 289 -1019
rect 89 -1069 289 -1053
rect 467 -1019 667 -972
rect 467 -1053 483 -1019
rect 651 -1053 667 -1019
rect 467 -1069 667 -1053
<< polycont >>
rect -651 1019 -483 1053
rect -273 1019 -105 1053
rect 105 1019 273 1053
rect 483 1019 651 1053
rect -651 691 -483 725
rect -273 691 -105 725
rect 105 691 273 725
rect 483 691 651 725
rect -651 583 -483 617
rect -273 583 -105 617
rect 105 583 273 617
rect 483 583 651 617
rect -651 255 -483 289
rect -273 255 -105 289
rect 105 255 273 289
rect 483 255 651 289
rect -651 147 -483 181
rect -273 147 -105 181
rect 105 147 273 181
rect 483 147 651 181
rect -651 -181 -483 -147
rect -273 -181 -105 -147
rect 105 -181 273 -147
rect 483 -181 651 -147
rect -651 -289 -483 -255
rect -273 -289 -105 -255
rect 105 -289 273 -255
rect 483 -289 651 -255
rect -651 -617 -483 -583
rect -273 -617 -105 -583
rect 105 -617 273 -583
rect 483 -617 651 -583
rect -651 -725 -483 -691
rect -273 -725 -105 -691
rect 105 -725 273 -691
rect 483 -725 651 -691
rect -651 -1053 -483 -1019
rect -273 -1053 -105 -1019
rect 105 -1053 273 -1019
rect 483 -1053 651 -1019
<< locali >>
rect -847 1157 -751 1191
rect 751 1157 847 1191
rect -847 1095 -813 1157
rect 813 1095 847 1157
rect -667 1019 -651 1053
rect -483 1019 -467 1053
rect -289 1019 -273 1053
rect -105 1019 -89 1053
rect 89 1019 105 1053
rect 273 1019 289 1053
rect 467 1019 483 1053
rect 651 1019 667 1053
rect -713 960 -679 976
rect -713 768 -679 784
rect -455 960 -421 976
rect -455 768 -421 784
rect -335 960 -301 976
rect -335 768 -301 784
rect -77 960 -43 976
rect -77 768 -43 784
rect 43 960 77 976
rect 43 768 77 784
rect 301 960 335 976
rect 301 768 335 784
rect 421 960 455 976
rect 421 768 455 784
rect 679 960 713 976
rect 679 768 713 784
rect -667 691 -651 725
rect -483 691 -467 725
rect -289 691 -273 725
rect -105 691 -89 725
rect 89 691 105 725
rect 273 691 289 725
rect 467 691 483 725
rect 651 691 667 725
rect -667 583 -651 617
rect -483 583 -467 617
rect -289 583 -273 617
rect -105 583 -89 617
rect 89 583 105 617
rect 273 583 289 617
rect 467 583 483 617
rect 651 583 667 617
rect -713 524 -679 540
rect -713 332 -679 348
rect -455 524 -421 540
rect -455 332 -421 348
rect -335 524 -301 540
rect -335 332 -301 348
rect -77 524 -43 540
rect -77 332 -43 348
rect 43 524 77 540
rect 43 332 77 348
rect 301 524 335 540
rect 301 332 335 348
rect 421 524 455 540
rect 421 332 455 348
rect 679 524 713 540
rect 679 332 713 348
rect -667 255 -651 289
rect -483 255 -467 289
rect -289 255 -273 289
rect -105 255 -89 289
rect 89 255 105 289
rect 273 255 289 289
rect 467 255 483 289
rect 651 255 667 289
rect -667 147 -651 181
rect -483 147 -467 181
rect -289 147 -273 181
rect -105 147 -89 181
rect 89 147 105 181
rect 273 147 289 181
rect 467 147 483 181
rect 651 147 667 181
rect -713 88 -679 104
rect -713 -104 -679 -88
rect -455 88 -421 104
rect -455 -104 -421 -88
rect -335 88 -301 104
rect -335 -104 -301 -88
rect -77 88 -43 104
rect -77 -104 -43 -88
rect 43 88 77 104
rect 43 -104 77 -88
rect 301 88 335 104
rect 301 -104 335 -88
rect 421 88 455 104
rect 421 -104 455 -88
rect 679 88 713 104
rect 679 -104 713 -88
rect -667 -181 -651 -147
rect -483 -181 -467 -147
rect -289 -181 -273 -147
rect -105 -181 -89 -147
rect 89 -181 105 -147
rect 273 -181 289 -147
rect 467 -181 483 -147
rect 651 -181 667 -147
rect -667 -289 -651 -255
rect -483 -289 -467 -255
rect -289 -289 -273 -255
rect -105 -289 -89 -255
rect 89 -289 105 -255
rect 273 -289 289 -255
rect 467 -289 483 -255
rect 651 -289 667 -255
rect -713 -348 -679 -332
rect -713 -540 -679 -524
rect -455 -348 -421 -332
rect -455 -540 -421 -524
rect -335 -348 -301 -332
rect -335 -540 -301 -524
rect -77 -348 -43 -332
rect -77 -540 -43 -524
rect 43 -348 77 -332
rect 43 -540 77 -524
rect 301 -348 335 -332
rect 301 -540 335 -524
rect 421 -348 455 -332
rect 421 -540 455 -524
rect 679 -348 713 -332
rect 679 -540 713 -524
rect -667 -617 -651 -583
rect -483 -617 -467 -583
rect -289 -617 -273 -583
rect -105 -617 -89 -583
rect 89 -617 105 -583
rect 273 -617 289 -583
rect 467 -617 483 -583
rect 651 -617 667 -583
rect -667 -725 -651 -691
rect -483 -725 -467 -691
rect -289 -725 -273 -691
rect -105 -725 -89 -691
rect 89 -725 105 -691
rect 273 -725 289 -691
rect 467 -725 483 -691
rect 651 -725 667 -691
rect -713 -784 -679 -768
rect -713 -976 -679 -960
rect -455 -784 -421 -768
rect -455 -976 -421 -960
rect -335 -784 -301 -768
rect -335 -976 -301 -960
rect -77 -784 -43 -768
rect -77 -976 -43 -960
rect 43 -784 77 -768
rect 43 -976 77 -960
rect 301 -784 335 -768
rect 301 -976 335 -960
rect 421 -784 455 -768
rect 421 -976 455 -960
rect 679 -784 713 -768
rect 679 -976 713 -960
rect -667 -1053 -651 -1019
rect -483 -1053 -467 -1019
rect -289 -1053 -273 -1019
rect -105 -1053 -89 -1019
rect 89 -1053 105 -1019
rect 273 -1053 289 -1019
rect 467 -1053 483 -1019
rect 651 -1053 667 -1019
rect -847 -1157 -813 -1095
rect 813 -1157 847 -1095
rect -847 -1191 -751 -1157
rect 751 -1191 847 -1157
<< viali >>
rect -651 1019 -483 1053
rect -273 1019 -105 1053
rect 105 1019 273 1053
rect 483 1019 651 1053
rect -713 784 -679 960
rect -455 784 -421 960
rect -335 784 -301 960
rect -77 784 -43 960
rect 43 784 77 960
rect 301 784 335 960
rect 421 784 455 960
rect 679 784 713 960
rect -651 691 -483 725
rect -273 691 -105 725
rect 105 691 273 725
rect 483 691 651 725
rect -651 583 -483 617
rect -273 583 -105 617
rect 105 583 273 617
rect 483 583 651 617
rect -713 348 -679 524
rect -455 348 -421 524
rect -335 348 -301 524
rect -77 348 -43 524
rect 43 348 77 524
rect 301 348 335 524
rect 421 348 455 524
rect 679 348 713 524
rect -651 255 -483 289
rect -273 255 -105 289
rect 105 255 273 289
rect 483 255 651 289
rect -651 147 -483 181
rect -273 147 -105 181
rect 105 147 273 181
rect 483 147 651 181
rect -713 -88 -679 88
rect -455 -88 -421 88
rect -335 -88 -301 88
rect -77 -88 -43 88
rect 43 -88 77 88
rect 301 -88 335 88
rect 421 -88 455 88
rect 679 -88 713 88
rect -651 -181 -483 -147
rect -273 -181 -105 -147
rect 105 -181 273 -147
rect 483 -181 651 -147
rect -651 -289 -483 -255
rect -273 -289 -105 -255
rect 105 -289 273 -255
rect 483 -289 651 -255
rect -713 -524 -679 -348
rect -455 -524 -421 -348
rect -335 -524 -301 -348
rect -77 -524 -43 -348
rect 43 -524 77 -348
rect 301 -524 335 -348
rect 421 -524 455 -348
rect 679 -524 713 -348
rect -651 -617 -483 -583
rect -273 -617 -105 -583
rect 105 -617 273 -583
rect 483 -617 651 -583
rect -651 -725 -483 -691
rect -273 -725 -105 -691
rect 105 -725 273 -691
rect 483 -725 651 -691
rect -713 -960 -679 -784
rect -455 -960 -421 -784
rect -335 -960 -301 -784
rect -77 -960 -43 -784
rect 43 -960 77 -784
rect 301 -960 335 -784
rect 421 -960 455 -784
rect 679 -960 713 -784
rect -651 -1053 -483 -1019
rect -273 -1053 -105 -1019
rect 105 -1053 273 -1019
rect 483 -1053 651 -1019
<< metal1 >>
rect -663 1053 -471 1059
rect -663 1019 -651 1053
rect -483 1019 -471 1053
rect -663 1013 -471 1019
rect -285 1053 -93 1059
rect -285 1019 -273 1053
rect -105 1019 -93 1053
rect -285 1013 -93 1019
rect 93 1053 285 1059
rect 93 1019 105 1053
rect 273 1019 285 1053
rect 93 1013 285 1019
rect 471 1053 663 1059
rect 471 1019 483 1053
rect 651 1019 663 1053
rect 471 1013 663 1019
rect -719 960 -673 972
rect -719 784 -713 960
rect -679 784 -673 960
rect -719 772 -673 784
rect -461 960 -415 972
rect -461 784 -455 960
rect -421 784 -415 960
rect -461 772 -415 784
rect -341 960 -295 972
rect -341 784 -335 960
rect -301 784 -295 960
rect -341 772 -295 784
rect -83 960 -37 972
rect -83 784 -77 960
rect -43 784 -37 960
rect -83 772 -37 784
rect 37 960 83 972
rect 37 784 43 960
rect 77 784 83 960
rect 37 772 83 784
rect 295 960 341 972
rect 295 784 301 960
rect 335 784 341 960
rect 295 772 341 784
rect 415 960 461 972
rect 415 784 421 960
rect 455 784 461 960
rect 415 772 461 784
rect 673 960 719 972
rect 673 784 679 960
rect 713 784 719 960
rect 673 772 719 784
rect -663 725 -471 731
rect -663 691 -651 725
rect -483 691 -471 725
rect -663 685 -471 691
rect -285 725 -93 731
rect -285 691 -273 725
rect -105 691 -93 725
rect -285 685 -93 691
rect 93 725 285 731
rect 93 691 105 725
rect 273 691 285 725
rect 93 685 285 691
rect 471 725 663 731
rect 471 691 483 725
rect 651 691 663 725
rect 471 685 663 691
rect -663 617 -471 623
rect -663 583 -651 617
rect -483 583 -471 617
rect -663 577 -471 583
rect -285 617 -93 623
rect -285 583 -273 617
rect -105 583 -93 617
rect -285 577 -93 583
rect 93 617 285 623
rect 93 583 105 617
rect 273 583 285 617
rect 93 577 285 583
rect 471 617 663 623
rect 471 583 483 617
rect 651 583 663 617
rect 471 577 663 583
rect -719 524 -673 536
rect -719 348 -713 524
rect -679 348 -673 524
rect -719 336 -673 348
rect -461 524 -415 536
rect -461 348 -455 524
rect -421 348 -415 524
rect -461 336 -415 348
rect -341 524 -295 536
rect -341 348 -335 524
rect -301 348 -295 524
rect -341 336 -295 348
rect -83 524 -37 536
rect -83 348 -77 524
rect -43 348 -37 524
rect -83 336 -37 348
rect 37 524 83 536
rect 37 348 43 524
rect 77 348 83 524
rect 37 336 83 348
rect 295 524 341 536
rect 295 348 301 524
rect 335 348 341 524
rect 295 336 341 348
rect 415 524 461 536
rect 415 348 421 524
rect 455 348 461 524
rect 415 336 461 348
rect 673 524 719 536
rect 673 348 679 524
rect 713 348 719 524
rect 673 336 719 348
rect -663 289 -471 295
rect -663 255 -651 289
rect -483 255 -471 289
rect -663 249 -471 255
rect -285 289 -93 295
rect -285 255 -273 289
rect -105 255 -93 289
rect -285 249 -93 255
rect 93 289 285 295
rect 93 255 105 289
rect 273 255 285 289
rect 93 249 285 255
rect 471 289 663 295
rect 471 255 483 289
rect 651 255 663 289
rect 471 249 663 255
rect -663 181 -471 187
rect -663 147 -651 181
rect -483 147 -471 181
rect -663 141 -471 147
rect -285 181 -93 187
rect -285 147 -273 181
rect -105 147 -93 181
rect -285 141 -93 147
rect 93 181 285 187
rect 93 147 105 181
rect 273 147 285 181
rect 93 141 285 147
rect 471 181 663 187
rect 471 147 483 181
rect 651 147 663 181
rect 471 141 663 147
rect -719 88 -673 100
rect -719 -88 -713 88
rect -679 -88 -673 88
rect -719 -100 -673 -88
rect -461 88 -415 100
rect -461 -88 -455 88
rect -421 -88 -415 88
rect -461 -100 -415 -88
rect -341 88 -295 100
rect -341 -88 -335 88
rect -301 -88 -295 88
rect -341 -100 -295 -88
rect -83 88 -37 100
rect -83 -88 -77 88
rect -43 -88 -37 88
rect -83 -100 -37 -88
rect 37 88 83 100
rect 37 -88 43 88
rect 77 -88 83 88
rect 37 -100 83 -88
rect 295 88 341 100
rect 295 -88 301 88
rect 335 -88 341 88
rect 295 -100 341 -88
rect 415 88 461 100
rect 415 -88 421 88
rect 455 -88 461 88
rect 415 -100 461 -88
rect 673 88 719 100
rect 673 -88 679 88
rect 713 -88 719 88
rect 673 -100 719 -88
rect -663 -147 -471 -141
rect -663 -181 -651 -147
rect -483 -181 -471 -147
rect -663 -187 -471 -181
rect -285 -147 -93 -141
rect -285 -181 -273 -147
rect -105 -181 -93 -147
rect -285 -187 -93 -181
rect 93 -147 285 -141
rect 93 -181 105 -147
rect 273 -181 285 -147
rect 93 -187 285 -181
rect 471 -147 663 -141
rect 471 -181 483 -147
rect 651 -181 663 -147
rect 471 -187 663 -181
rect -663 -255 -471 -249
rect -663 -289 -651 -255
rect -483 -289 -471 -255
rect -663 -295 -471 -289
rect -285 -255 -93 -249
rect -285 -289 -273 -255
rect -105 -289 -93 -255
rect -285 -295 -93 -289
rect 93 -255 285 -249
rect 93 -289 105 -255
rect 273 -289 285 -255
rect 93 -295 285 -289
rect 471 -255 663 -249
rect 471 -289 483 -255
rect 651 -289 663 -255
rect 471 -295 663 -289
rect -719 -348 -673 -336
rect -719 -524 -713 -348
rect -679 -524 -673 -348
rect -719 -536 -673 -524
rect -461 -348 -415 -336
rect -461 -524 -455 -348
rect -421 -524 -415 -348
rect -461 -536 -415 -524
rect -341 -348 -295 -336
rect -341 -524 -335 -348
rect -301 -524 -295 -348
rect -341 -536 -295 -524
rect -83 -348 -37 -336
rect -83 -524 -77 -348
rect -43 -524 -37 -348
rect -83 -536 -37 -524
rect 37 -348 83 -336
rect 37 -524 43 -348
rect 77 -524 83 -348
rect 37 -536 83 -524
rect 295 -348 341 -336
rect 295 -524 301 -348
rect 335 -524 341 -348
rect 295 -536 341 -524
rect 415 -348 461 -336
rect 415 -524 421 -348
rect 455 -524 461 -348
rect 415 -536 461 -524
rect 673 -348 719 -336
rect 673 -524 679 -348
rect 713 -524 719 -348
rect 673 -536 719 -524
rect -663 -583 -471 -577
rect -663 -617 -651 -583
rect -483 -617 -471 -583
rect -663 -623 -471 -617
rect -285 -583 -93 -577
rect -285 -617 -273 -583
rect -105 -617 -93 -583
rect -285 -623 -93 -617
rect 93 -583 285 -577
rect 93 -617 105 -583
rect 273 -617 285 -583
rect 93 -623 285 -617
rect 471 -583 663 -577
rect 471 -617 483 -583
rect 651 -617 663 -583
rect 471 -623 663 -617
rect -663 -691 -471 -685
rect -663 -725 -651 -691
rect -483 -725 -471 -691
rect -663 -731 -471 -725
rect -285 -691 -93 -685
rect -285 -725 -273 -691
rect -105 -725 -93 -691
rect -285 -731 -93 -725
rect 93 -691 285 -685
rect 93 -725 105 -691
rect 273 -725 285 -691
rect 93 -731 285 -725
rect 471 -691 663 -685
rect 471 -725 483 -691
rect 651 -725 663 -691
rect 471 -731 663 -725
rect -719 -784 -673 -772
rect -719 -960 -713 -784
rect -679 -960 -673 -784
rect -719 -972 -673 -960
rect -461 -784 -415 -772
rect -461 -960 -455 -784
rect -421 -960 -415 -784
rect -461 -972 -415 -960
rect -341 -784 -295 -772
rect -341 -960 -335 -784
rect -301 -960 -295 -784
rect -341 -972 -295 -960
rect -83 -784 -37 -772
rect -83 -960 -77 -784
rect -43 -960 -37 -784
rect -83 -972 -37 -960
rect 37 -784 83 -772
rect 37 -960 43 -784
rect 77 -960 83 -784
rect 37 -972 83 -960
rect 295 -784 341 -772
rect 295 -960 301 -784
rect 335 -960 341 -784
rect 295 -972 341 -960
rect 415 -784 461 -772
rect 415 -960 421 -784
rect 455 -960 461 -784
rect 415 -972 461 -960
rect 673 -784 719 -772
rect 673 -960 679 -784
rect 713 -960 719 -784
rect 673 -972 719 -960
rect -663 -1019 -471 -1013
rect -663 -1053 -651 -1019
rect -483 -1053 -471 -1019
rect -663 -1059 -471 -1053
rect -285 -1019 -93 -1013
rect -285 -1053 -273 -1019
rect -105 -1053 -93 -1019
rect -285 -1059 -93 -1053
rect 93 -1019 285 -1013
rect 93 -1053 105 -1019
rect 273 -1053 285 -1019
rect 93 -1059 285 -1053
rect 471 -1019 663 -1013
rect 471 -1053 483 -1019
rect 651 -1053 663 -1019
rect 471 -1059 663 -1053
<< properties >>
string FIXED_BBOX -830 -1174 830 1174
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
