magic
tech sky130A
magscale 1 2
timestamp 1628260645
<< pwell >>
rect -201 -1598 201 1598
<< psubdiff >>
rect -165 1528 -69 1562
rect 69 1528 165 1562
rect -165 1466 -131 1528
rect 131 1466 165 1528
rect -165 -1528 -131 -1466
rect 131 -1528 165 -1466
rect -165 -1562 -69 -1528
rect 69 -1562 165 -1528
<< psubdiffcont >>
rect -69 1528 69 1562
rect -165 -1466 -131 1466
rect 131 -1466 165 1466
rect -69 -1562 69 -1528
<< xpolycontact >>
rect -35 1000 35 1432
rect -35 -1432 35 -1000
<< xpolyres >>
rect -35 -1000 35 1000
<< locali >>
rect -165 1528 -69 1562
rect 69 1528 165 1562
rect -165 1466 -131 1528
rect 131 1466 165 1528
rect -165 -1528 -131 -1466
rect 131 -1528 165 -1466
rect -165 -1562 -69 -1528
rect 69 -1562 165 -1528
<< viali >>
rect -19 1017 19 1414
rect -19 -1414 19 -1017
<< metal1 >>
rect -25 1414 25 1426
rect -25 1017 -19 1414
rect 19 1017 25 1414
rect -25 1005 25 1017
rect -25 -1017 25 -1005
rect -25 -1414 -19 -1017
rect 19 -1414 25 -1017
rect -25 -1426 25 -1414
<< res0p35 >>
rect -37 -1002 37 1002
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string FIXED_BBOX -148 -1545 148 1545
string parameters w 0.350 l 10 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 57.252k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
