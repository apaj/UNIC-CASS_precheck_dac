* NGSPICE file created from dac_cell1.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p69_MS44J6 a_n69_n6232# a_n69_5800# a_n199_n6362#
X0 a_n69_5800# a_n69_n6232# a_n199_n6362# sky130_fd_pr__res_xhigh_po_0p69 l=58
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0 a_n100_n197# a_100_n100# w_n358_n397#
+ a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n358_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt dac_cell1 vsup vgnd iref vsw iout iout_n vbias
XXR1 parR sourceM2 vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXR2 parR sourceM2 vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXR4 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0
XXM2 iref sourceM3M4 vsup sourceM2 sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0
XXM3 vsw iout vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0
XXM4 vbias iout_n vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0
.ends

