magic
tech sky130A
timestamp 1628499526
<< pwell >>
rect -139 -2529 139 2529
<< mvnmos >>
rect -25 -2400 25 2400
<< mvndiff >>
rect -54 2394 -25 2400
rect -54 -2394 -48 2394
rect -31 -2394 -25 2394
rect -54 -2400 -25 -2394
rect 25 2394 54 2400
rect 25 -2394 31 2394
rect 48 -2394 54 2394
rect 25 -2400 54 -2394
<< mvndiffc >>
rect -48 -2394 -31 2394
rect 31 -2394 48 2394
<< mvpsubdiff >>
rect -121 2505 121 2511
rect -121 2488 -67 2505
rect 67 2488 121 2505
rect -121 2482 121 2488
rect -121 2457 -92 2482
rect -121 -2457 -115 2457
rect -98 -2457 -92 2457
rect 92 2457 121 2482
rect -121 -2482 -92 -2457
rect 92 -2457 98 2457
rect 115 -2457 121 2457
rect 92 -2482 121 -2457
rect -121 -2488 121 -2482
rect -121 -2505 -67 -2488
rect 67 -2505 121 -2488
rect -121 -2511 121 -2505
<< mvpsubdiffcont >>
rect -67 2488 67 2505
rect -115 -2457 -98 2457
rect 98 -2457 115 2457
rect -67 -2505 67 -2488
<< poly >>
rect -25 2436 25 2444
rect -25 2419 -17 2436
rect 17 2419 25 2436
rect -25 2400 25 2419
rect -25 -2419 25 -2400
rect -25 -2436 -17 -2419
rect 17 -2436 25 -2419
rect -25 -2444 25 -2436
<< polycont >>
rect -17 2419 17 2436
rect -17 -2436 17 -2419
<< locali >>
rect -115 2488 -67 2505
rect 67 2488 115 2505
rect -115 2457 -98 2488
rect 98 2457 115 2488
rect -25 2419 -17 2436
rect 17 2419 25 2436
rect -48 2394 -31 2402
rect -48 -2402 -31 -2394
rect 31 2394 48 2402
rect 31 -2402 48 -2394
rect -25 -2436 -17 -2419
rect 17 -2436 25 -2419
rect -115 -2488 -98 -2457
rect 98 -2488 115 -2457
rect -115 -2505 -67 -2488
rect 67 -2505 115 -2488
<< viali >>
rect -17 2419 17 2436
rect -48 -2394 -31 2394
rect 31 -2394 48 2394
rect -17 -2436 17 -2419
<< metal1 >>
rect -23 2436 23 2439
rect -23 2419 -17 2436
rect 17 2419 23 2436
rect -23 2416 23 2419
rect -51 2394 -28 2400
rect -51 -2394 -48 2394
rect -31 -2394 -28 2394
rect -51 -2400 -28 -2394
rect 28 2394 51 2400
rect 28 -2394 31 2394
rect 48 -2394 51 2394
rect 28 -2400 51 -2394
rect -23 -2419 23 -2416
rect -23 -2436 -17 -2419
rect 17 -2436 23 -2419
rect -23 -2439 23 -2436
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -106 -2496 106 2496
string parameters w 48 l 0.50 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
