* SPICE3 file created from dac_cell4.ext - technology: sky130A

.option scale=5000u

.subckt dac_cell4 vsup vgnd iref vsw iout iout_n vbias
X0 m1_3264_4148# li_984_4388# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=1260
X1 m1_3264_4148# li_984_4388# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=1260
X2 m1_3264_4148# vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=1260
X3 m1_3264_4148# vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=1260
X4 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 ad=11600 pd=516 as=290000 ps=10464 w=200 l=200
X5 vsup iref li_984_4388# vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1600 l=200
X6 iout vsw vsup vsup sky130_fd_pr__pfet_g5v0d10v5 ad=92800 pd=3316 as=0 ps=0 w=1600 l=200
X7 iout_n vbias vsup vsup sky130_fd_pr__pfet_g5v0d10v5 ad=92800 pd=3316 as=0 ps=0 w=1600 l=200
.ends
