magic
tech sky130A
magscale 1 2
timestamp 1696881349
<< nwell >>
rect -925 -1051 925 1051
<< mvpmos >>
rect -667 554 -467 754
rect -289 554 -89 754
rect 89 554 289 754
rect 467 554 667 754
rect -667 118 -467 318
rect -289 118 -89 318
rect 89 118 289 318
rect 467 118 667 318
rect -667 -318 -467 -118
rect -289 -318 -89 -118
rect 89 -318 289 -118
rect 467 -318 667 -118
rect -667 -754 -467 -554
rect -289 -754 -89 -554
rect 89 -754 289 -554
rect 467 -754 667 -554
<< mvpdiff >>
rect -725 742 -667 754
rect -725 566 -713 742
rect -679 566 -667 742
rect -725 554 -667 566
rect -467 742 -409 754
rect -467 566 -455 742
rect -421 566 -409 742
rect -467 554 -409 566
rect -347 742 -289 754
rect -347 566 -335 742
rect -301 566 -289 742
rect -347 554 -289 566
rect -89 742 -31 754
rect -89 566 -77 742
rect -43 566 -31 742
rect -89 554 -31 566
rect 31 742 89 754
rect 31 566 43 742
rect 77 566 89 742
rect 31 554 89 566
rect 289 742 347 754
rect 289 566 301 742
rect 335 566 347 742
rect 289 554 347 566
rect 409 742 467 754
rect 409 566 421 742
rect 455 566 467 742
rect 409 554 467 566
rect 667 742 725 754
rect 667 566 679 742
rect 713 566 725 742
rect 667 554 725 566
rect -725 306 -667 318
rect -725 130 -713 306
rect -679 130 -667 306
rect -725 118 -667 130
rect -467 306 -409 318
rect -467 130 -455 306
rect -421 130 -409 306
rect -467 118 -409 130
rect -347 306 -289 318
rect -347 130 -335 306
rect -301 130 -289 306
rect -347 118 -289 130
rect -89 306 -31 318
rect -89 130 -77 306
rect -43 130 -31 306
rect -89 118 -31 130
rect 31 306 89 318
rect 31 130 43 306
rect 77 130 89 306
rect 31 118 89 130
rect 289 306 347 318
rect 289 130 301 306
rect 335 130 347 306
rect 289 118 347 130
rect 409 306 467 318
rect 409 130 421 306
rect 455 130 467 306
rect 409 118 467 130
rect 667 306 725 318
rect 667 130 679 306
rect 713 130 725 306
rect 667 118 725 130
rect -725 -130 -667 -118
rect -725 -306 -713 -130
rect -679 -306 -667 -130
rect -725 -318 -667 -306
rect -467 -130 -409 -118
rect -467 -306 -455 -130
rect -421 -306 -409 -130
rect -467 -318 -409 -306
rect -347 -130 -289 -118
rect -347 -306 -335 -130
rect -301 -306 -289 -130
rect -347 -318 -289 -306
rect -89 -130 -31 -118
rect -89 -306 -77 -130
rect -43 -306 -31 -130
rect -89 -318 -31 -306
rect 31 -130 89 -118
rect 31 -306 43 -130
rect 77 -306 89 -130
rect 31 -318 89 -306
rect 289 -130 347 -118
rect 289 -306 301 -130
rect 335 -306 347 -130
rect 289 -318 347 -306
rect 409 -130 467 -118
rect 409 -306 421 -130
rect 455 -306 467 -130
rect 409 -318 467 -306
rect 667 -130 725 -118
rect 667 -306 679 -130
rect 713 -306 725 -130
rect 667 -318 725 -306
rect -725 -566 -667 -554
rect -725 -742 -713 -566
rect -679 -742 -667 -566
rect -725 -754 -667 -742
rect -467 -566 -409 -554
rect -467 -742 -455 -566
rect -421 -742 -409 -566
rect -467 -754 -409 -742
rect -347 -566 -289 -554
rect -347 -742 -335 -566
rect -301 -742 -289 -566
rect -347 -754 -289 -742
rect -89 -566 -31 -554
rect -89 -742 -77 -566
rect -43 -742 -31 -566
rect -89 -754 -31 -742
rect 31 -566 89 -554
rect 31 -742 43 -566
rect 77 -742 89 -566
rect 31 -754 89 -742
rect 289 -566 347 -554
rect 289 -742 301 -566
rect 335 -742 347 -566
rect 289 -754 347 -742
rect 409 -566 467 -554
rect 409 -742 421 -566
rect 455 -742 467 -566
rect 409 -754 467 -742
rect 667 -566 725 -554
rect 667 -742 679 -566
rect 713 -742 725 -566
rect 667 -754 725 -742
<< mvpdiffc >>
rect -713 566 -679 742
rect -455 566 -421 742
rect -335 566 -301 742
rect -77 566 -43 742
rect 43 566 77 742
rect 301 566 335 742
rect 421 566 455 742
rect 679 566 713 742
rect -713 130 -679 306
rect -455 130 -421 306
rect -335 130 -301 306
rect -77 130 -43 306
rect 43 130 77 306
rect 301 130 335 306
rect 421 130 455 306
rect 679 130 713 306
rect -713 -306 -679 -130
rect -455 -306 -421 -130
rect -335 -306 -301 -130
rect -77 -306 -43 -130
rect 43 -306 77 -130
rect 301 -306 335 -130
rect 421 -306 455 -130
rect 679 -306 713 -130
rect -713 -742 -679 -566
rect -455 -742 -421 -566
rect -335 -742 -301 -566
rect -77 -742 -43 -566
rect 43 -742 77 -566
rect 301 -742 335 -566
rect 421 -742 455 -566
rect 679 -742 713 -566
<< mvnsubdiff >>
rect -859 973 859 985
rect -859 939 -751 973
rect 751 939 859 973
rect -859 927 859 939
rect -859 877 -801 927
rect -859 -877 -847 877
rect -813 -877 -801 877
rect 801 877 859 927
rect -859 -927 -801 -877
rect 801 -877 813 877
rect 847 -877 859 877
rect 801 -927 859 -877
rect -859 -939 859 -927
rect -859 -973 -751 -939
rect 751 -973 859 -939
rect -859 -985 859 -973
<< mvnsubdiffcont >>
rect -751 939 751 973
rect -847 -877 -813 877
rect 813 -877 847 877
rect -751 -973 751 -939
<< poly >>
rect -667 835 -467 851
rect -667 801 -651 835
rect -483 801 -467 835
rect -667 754 -467 801
rect -289 835 -89 851
rect -289 801 -273 835
rect -105 801 -89 835
rect -289 754 -89 801
rect 89 835 289 851
rect 89 801 105 835
rect 273 801 289 835
rect 89 754 289 801
rect 467 835 667 851
rect 467 801 483 835
rect 651 801 667 835
rect 467 754 667 801
rect -667 507 -467 554
rect -667 473 -651 507
rect -483 473 -467 507
rect -667 457 -467 473
rect -289 507 -89 554
rect -289 473 -273 507
rect -105 473 -89 507
rect -289 457 -89 473
rect 89 507 289 554
rect 89 473 105 507
rect 273 473 289 507
rect 89 457 289 473
rect 467 507 667 554
rect 467 473 483 507
rect 651 473 667 507
rect 467 457 667 473
rect -667 399 -467 415
rect -667 365 -651 399
rect -483 365 -467 399
rect -667 318 -467 365
rect -289 399 -89 415
rect -289 365 -273 399
rect -105 365 -89 399
rect -289 318 -89 365
rect 89 399 289 415
rect 89 365 105 399
rect 273 365 289 399
rect 89 318 289 365
rect 467 399 667 415
rect 467 365 483 399
rect 651 365 667 399
rect 467 318 667 365
rect -667 71 -467 118
rect -667 37 -651 71
rect -483 37 -467 71
rect -667 21 -467 37
rect -289 71 -89 118
rect -289 37 -273 71
rect -105 37 -89 71
rect -289 21 -89 37
rect 89 71 289 118
rect 89 37 105 71
rect 273 37 289 71
rect 89 21 289 37
rect 467 71 667 118
rect 467 37 483 71
rect 651 37 667 71
rect 467 21 667 37
rect -667 -37 -467 -21
rect -667 -71 -651 -37
rect -483 -71 -467 -37
rect -667 -118 -467 -71
rect -289 -37 -89 -21
rect -289 -71 -273 -37
rect -105 -71 -89 -37
rect -289 -118 -89 -71
rect 89 -37 289 -21
rect 89 -71 105 -37
rect 273 -71 289 -37
rect 89 -118 289 -71
rect 467 -37 667 -21
rect 467 -71 483 -37
rect 651 -71 667 -37
rect 467 -118 667 -71
rect -667 -365 -467 -318
rect -667 -399 -651 -365
rect -483 -399 -467 -365
rect -667 -415 -467 -399
rect -289 -365 -89 -318
rect -289 -399 -273 -365
rect -105 -399 -89 -365
rect -289 -415 -89 -399
rect 89 -365 289 -318
rect 89 -399 105 -365
rect 273 -399 289 -365
rect 89 -415 289 -399
rect 467 -365 667 -318
rect 467 -399 483 -365
rect 651 -399 667 -365
rect 467 -415 667 -399
rect -667 -473 -467 -457
rect -667 -507 -651 -473
rect -483 -507 -467 -473
rect -667 -554 -467 -507
rect -289 -473 -89 -457
rect -289 -507 -273 -473
rect -105 -507 -89 -473
rect -289 -554 -89 -507
rect 89 -473 289 -457
rect 89 -507 105 -473
rect 273 -507 289 -473
rect 89 -554 289 -507
rect 467 -473 667 -457
rect 467 -507 483 -473
rect 651 -507 667 -473
rect 467 -554 667 -507
rect -667 -801 -467 -754
rect -667 -835 -651 -801
rect -483 -835 -467 -801
rect -667 -851 -467 -835
rect -289 -801 -89 -754
rect -289 -835 -273 -801
rect -105 -835 -89 -801
rect -289 -851 -89 -835
rect 89 -801 289 -754
rect 89 -835 105 -801
rect 273 -835 289 -801
rect 89 -851 289 -835
rect 467 -801 667 -754
rect 467 -835 483 -801
rect 651 -835 667 -801
rect 467 -851 667 -835
<< polycont >>
rect -651 801 -483 835
rect -273 801 -105 835
rect 105 801 273 835
rect 483 801 651 835
rect -651 473 -483 507
rect -273 473 -105 507
rect 105 473 273 507
rect 483 473 651 507
rect -651 365 -483 399
rect -273 365 -105 399
rect 105 365 273 399
rect 483 365 651 399
rect -651 37 -483 71
rect -273 37 -105 71
rect 105 37 273 71
rect 483 37 651 71
rect -651 -71 -483 -37
rect -273 -71 -105 -37
rect 105 -71 273 -37
rect 483 -71 651 -37
rect -651 -399 -483 -365
rect -273 -399 -105 -365
rect 105 -399 273 -365
rect 483 -399 651 -365
rect -651 -507 -483 -473
rect -273 -507 -105 -473
rect 105 -507 273 -473
rect 483 -507 651 -473
rect -651 -835 -483 -801
rect -273 -835 -105 -801
rect 105 -835 273 -801
rect 483 -835 651 -801
<< locali >>
rect -847 939 -751 973
rect 751 939 847 973
rect -847 877 -813 939
rect 813 877 847 939
rect -667 801 -651 835
rect -483 801 -467 835
rect -289 801 -273 835
rect -105 801 -89 835
rect 89 801 105 835
rect 273 801 289 835
rect 467 801 483 835
rect 651 801 667 835
rect -713 742 -679 758
rect -713 550 -679 566
rect -455 742 -421 758
rect -455 550 -421 566
rect -335 742 -301 758
rect -335 550 -301 566
rect -77 742 -43 758
rect -77 550 -43 566
rect 43 742 77 758
rect 43 550 77 566
rect 301 742 335 758
rect 301 550 335 566
rect 421 742 455 758
rect 421 550 455 566
rect 679 742 713 758
rect 679 550 713 566
rect -667 473 -651 507
rect -483 473 -467 507
rect -289 473 -273 507
rect -105 473 -89 507
rect 89 473 105 507
rect 273 473 289 507
rect 467 473 483 507
rect 651 473 667 507
rect -667 365 -651 399
rect -483 365 -467 399
rect -289 365 -273 399
rect -105 365 -89 399
rect 89 365 105 399
rect 273 365 289 399
rect 467 365 483 399
rect 651 365 667 399
rect -713 306 -679 322
rect -713 114 -679 130
rect -455 306 -421 322
rect -455 114 -421 130
rect -335 306 -301 322
rect -335 114 -301 130
rect -77 306 -43 322
rect -77 114 -43 130
rect 43 306 77 322
rect 43 114 77 130
rect 301 306 335 322
rect 301 114 335 130
rect 421 306 455 322
rect 421 114 455 130
rect 679 306 713 322
rect 679 114 713 130
rect -667 37 -651 71
rect -483 37 -467 71
rect -289 37 -273 71
rect -105 37 -89 71
rect 89 37 105 71
rect 273 37 289 71
rect 467 37 483 71
rect 651 37 667 71
rect -667 -71 -651 -37
rect -483 -71 -467 -37
rect -289 -71 -273 -37
rect -105 -71 -89 -37
rect 89 -71 105 -37
rect 273 -71 289 -37
rect 467 -71 483 -37
rect 651 -71 667 -37
rect -713 -130 -679 -114
rect -713 -322 -679 -306
rect -455 -130 -421 -114
rect -455 -322 -421 -306
rect -335 -130 -301 -114
rect -335 -322 -301 -306
rect -77 -130 -43 -114
rect -77 -322 -43 -306
rect 43 -130 77 -114
rect 43 -322 77 -306
rect 301 -130 335 -114
rect 301 -322 335 -306
rect 421 -130 455 -114
rect 421 -322 455 -306
rect 679 -130 713 -114
rect 679 -322 713 -306
rect -667 -399 -651 -365
rect -483 -399 -467 -365
rect -289 -399 -273 -365
rect -105 -399 -89 -365
rect 89 -399 105 -365
rect 273 -399 289 -365
rect 467 -399 483 -365
rect 651 -399 667 -365
rect -667 -507 -651 -473
rect -483 -507 -467 -473
rect -289 -507 -273 -473
rect -105 -507 -89 -473
rect 89 -507 105 -473
rect 273 -507 289 -473
rect 467 -507 483 -473
rect 651 -507 667 -473
rect -713 -566 -679 -550
rect -713 -758 -679 -742
rect -455 -566 -421 -550
rect -455 -758 -421 -742
rect -335 -566 -301 -550
rect -335 -758 -301 -742
rect -77 -566 -43 -550
rect -77 -758 -43 -742
rect 43 -566 77 -550
rect 43 -758 77 -742
rect 301 -566 335 -550
rect 301 -758 335 -742
rect 421 -566 455 -550
rect 421 -758 455 -742
rect 679 -566 713 -550
rect 679 -758 713 -742
rect -667 -835 -651 -801
rect -483 -835 -467 -801
rect -289 -835 -273 -801
rect -105 -835 -89 -801
rect 89 -835 105 -801
rect 273 -835 289 -801
rect 467 -835 483 -801
rect 651 -835 667 -801
rect -847 -939 -813 -877
rect 813 -939 847 -877
rect -847 -973 -751 -939
rect 751 -973 847 -939
<< viali >>
rect -651 801 -483 835
rect -273 801 -105 835
rect 105 801 273 835
rect 483 801 651 835
rect -713 566 -679 742
rect -455 566 -421 742
rect -335 566 -301 742
rect -77 566 -43 742
rect 43 566 77 742
rect 301 566 335 742
rect 421 566 455 742
rect 679 566 713 742
rect -651 473 -483 507
rect -273 473 -105 507
rect 105 473 273 507
rect 483 473 651 507
rect -651 365 -483 399
rect -273 365 -105 399
rect 105 365 273 399
rect 483 365 651 399
rect -713 130 -679 306
rect -455 130 -421 306
rect -335 130 -301 306
rect -77 130 -43 306
rect 43 130 77 306
rect 301 130 335 306
rect 421 130 455 306
rect 679 130 713 306
rect -651 37 -483 71
rect -273 37 -105 71
rect 105 37 273 71
rect 483 37 651 71
rect -651 -71 -483 -37
rect -273 -71 -105 -37
rect 105 -71 273 -37
rect 483 -71 651 -37
rect -713 -306 -679 -130
rect -455 -306 -421 -130
rect -335 -306 -301 -130
rect -77 -306 -43 -130
rect 43 -306 77 -130
rect 301 -306 335 -130
rect 421 -306 455 -130
rect 679 -306 713 -130
rect -651 -399 -483 -365
rect -273 -399 -105 -365
rect 105 -399 273 -365
rect 483 -399 651 -365
rect -651 -507 -483 -473
rect -273 -507 -105 -473
rect 105 -507 273 -473
rect 483 -507 651 -473
rect -713 -742 -679 -566
rect -455 -742 -421 -566
rect -335 -742 -301 -566
rect -77 -742 -43 -566
rect 43 -742 77 -566
rect 301 -742 335 -566
rect 421 -742 455 -566
rect 679 -742 713 -566
rect -651 -835 -483 -801
rect -273 -835 -105 -801
rect 105 -835 273 -801
rect 483 -835 651 -801
<< metal1 >>
rect -663 835 -471 841
rect -663 801 -651 835
rect -483 801 -471 835
rect -663 795 -471 801
rect -285 835 -93 841
rect -285 801 -273 835
rect -105 801 -93 835
rect -285 795 -93 801
rect 93 835 285 841
rect 93 801 105 835
rect 273 801 285 835
rect 93 795 285 801
rect 471 835 663 841
rect 471 801 483 835
rect 651 801 663 835
rect 471 795 663 801
rect -719 742 -673 754
rect -719 566 -713 742
rect -679 566 -673 742
rect -719 554 -673 566
rect -461 742 -415 754
rect -461 566 -455 742
rect -421 566 -415 742
rect -461 554 -415 566
rect -341 742 -295 754
rect -341 566 -335 742
rect -301 566 -295 742
rect -341 554 -295 566
rect -83 742 -37 754
rect -83 566 -77 742
rect -43 566 -37 742
rect -83 554 -37 566
rect 37 742 83 754
rect 37 566 43 742
rect 77 566 83 742
rect 37 554 83 566
rect 295 742 341 754
rect 295 566 301 742
rect 335 566 341 742
rect 295 554 341 566
rect 415 742 461 754
rect 415 566 421 742
rect 455 566 461 742
rect 415 554 461 566
rect 673 742 719 754
rect 673 566 679 742
rect 713 566 719 742
rect 673 554 719 566
rect -663 507 -471 513
rect -663 473 -651 507
rect -483 473 -471 507
rect -663 467 -471 473
rect -285 507 -93 513
rect -285 473 -273 507
rect -105 473 -93 507
rect -285 467 -93 473
rect 93 507 285 513
rect 93 473 105 507
rect 273 473 285 507
rect 93 467 285 473
rect 471 507 663 513
rect 471 473 483 507
rect 651 473 663 507
rect 471 467 663 473
rect -663 399 -471 405
rect -663 365 -651 399
rect -483 365 -471 399
rect -663 359 -471 365
rect -285 399 -93 405
rect -285 365 -273 399
rect -105 365 -93 399
rect -285 359 -93 365
rect 93 399 285 405
rect 93 365 105 399
rect 273 365 285 399
rect 93 359 285 365
rect 471 399 663 405
rect 471 365 483 399
rect 651 365 663 399
rect 471 359 663 365
rect -719 306 -673 318
rect -719 130 -713 306
rect -679 130 -673 306
rect -719 118 -673 130
rect -461 306 -415 318
rect -461 130 -455 306
rect -421 130 -415 306
rect -461 118 -415 130
rect -341 306 -295 318
rect -341 130 -335 306
rect -301 130 -295 306
rect -341 118 -295 130
rect -83 306 -37 318
rect -83 130 -77 306
rect -43 130 -37 306
rect -83 118 -37 130
rect 37 306 83 318
rect 37 130 43 306
rect 77 130 83 306
rect 37 118 83 130
rect 295 306 341 318
rect 295 130 301 306
rect 335 130 341 306
rect 295 118 341 130
rect 415 306 461 318
rect 415 130 421 306
rect 455 130 461 306
rect 415 118 461 130
rect 673 306 719 318
rect 673 130 679 306
rect 713 130 719 306
rect 673 118 719 130
rect -663 71 -471 77
rect -663 37 -651 71
rect -483 37 -471 71
rect -663 31 -471 37
rect -285 71 -93 77
rect -285 37 -273 71
rect -105 37 -93 71
rect -285 31 -93 37
rect 93 71 285 77
rect 93 37 105 71
rect 273 37 285 71
rect 93 31 285 37
rect 471 71 663 77
rect 471 37 483 71
rect 651 37 663 71
rect 471 31 663 37
rect -663 -37 -471 -31
rect -663 -71 -651 -37
rect -483 -71 -471 -37
rect -663 -77 -471 -71
rect -285 -37 -93 -31
rect -285 -71 -273 -37
rect -105 -71 -93 -37
rect -285 -77 -93 -71
rect 93 -37 285 -31
rect 93 -71 105 -37
rect 273 -71 285 -37
rect 93 -77 285 -71
rect 471 -37 663 -31
rect 471 -71 483 -37
rect 651 -71 663 -37
rect 471 -77 663 -71
rect -719 -130 -673 -118
rect -719 -306 -713 -130
rect -679 -306 -673 -130
rect -719 -318 -673 -306
rect -461 -130 -415 -118
rect -461 -306 -455 -130
rect -421 -306 -415 -130
rect -461 -318 -415 -306
rect -341 -130 -295 -118
rect -341 -306 -335 -130
rect -301 -306 -295 -130
rect -341 -318 -295 -306
rect -83 -130 -37 -118
rect -83 -306 -77 -130
rect -43 -306 -37 -130
rect -83 -318 -37 -306
rect 37 -130 83 -118
rect 37 -306 43 -130
rect 77 -306 83 -130
rect 37 -318 83 -306
rect 295 -130 341 -118
rect 295 -306 301 -130
rect 335 -306 341 -130
rect 295 -318 341 -306
rect 415 -130 461 -118
rect 415 -306 421 -130
rect 455 -306 461 -130
rect 415 -318 461 -306
rect 673 -130 719 -118
rect 673 -306 679 -130
rect 713 -306 719 -130
rect 673 -318 719 -306
rect -663 -365 -471 -359
rect -663 -399 -651 -365
rect -483 -399 -471 -365
rect -663 -405 -471 -399
rect -285 -365 -93 -359
rect -285 -399 -273 -365
rect -105 -399 -93 -365
rect -285 -405 -93 -399
rect 93 -365 285 -359
rect 93 -399 105 -365
rect 273 -399 285 -365
rect 93 -405 285 -399
rect 471 -365 663 -359
rect 471 -399 483 -365
rect 651 -399 663 -365
rect 471 -405 663 -399
rect -663 -473 -471 -467
rect -663 -507 -651 -473
rect -483 -507 -471 -473
rect -663 -513 -471 -507
rect -285 -473 -93 -467
rect -285 -507 -273 -473
rect -105 -507 -93 -473
rect -285 -513 -93 -507
rect 93 -473 285 -467
rect 93 -507 105 -473
rect 273 -507 285 -473
rect 93 -513 285 -507
rect 471 -473 663 -467
rect 471 -507 483 -473
rect 651 -507 663 -473
rect 471 -513 663 -507
rect -719 -566 -673 -554
rect -719 -742 -713 -566
rect -679 -742 -673 -566
rect -719 -754 -673 -742
rect -461 -566 -415 -554
rect -461 -742 -455 -566
rect -421 -742 -415 -566
rect -461 -754 -415 -742
rect -341 -566 -295 -554
rect -341 -742 -335 -566
rect -301 -742 -295 -566
rect -341 -754 -295 -742
rect -83 -566 -37 -554
rect -83 -742 -77 -566
rect -43 -742 -37 -566
rect -83 -754 -37 -742
rect 37 -566 83 -554
rect 37 -742 43 -566
rect 77 -742 83 -566
rect 37 -754 83 -742
rect 295 -566 341 -554
rect 295 -742 301 -566
rect 335 -742 341 -566
rect 295 -754 341 -742
rect 415 -566 461 -554
rect 415 -742 421 -566
rect 455 -742 461 -566
rect 415 -754 461 -742
rect 673 -566 719 -554
rect 673 -742 679 -566
rect 713 -742 719 -566
rect 673 -754 719 -742
rect -663 -801 -471 -795
rect -663 -835 -651 -801
rect -483 -835 -471 -801
rect -663 -841 -471 -835
rect -285 -801 -93 -795
rect -285 -835 -273 -801
rect -105 -835 -93 -801
rect -285 -841 -93 -835
rect 93 -801 285 -795
rect 93 -835 105 -801
rect 273 -835 285 -801
rect 93 -841 285 -835
rect 471 -801 663 -795
rect 471 -835 483 -801
rect 651 -835 663 -801
rect 471 -841 663 -835
<< properties >>
string FIXED_BBOX -830 -956 830 956
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 4 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
