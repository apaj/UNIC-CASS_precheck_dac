magic
tech sky130A
magscale 1 2
timestamp 1628235594
<< pwell >>
rect -692 -1367 692 1367
<< nnmos >>
rect -464 109 -364 1109
rect -188 109 -88 1109
rect 88 109 188 1109
rect 364 109 464 1109
rect -464 -1109 -364 -109
rect -188 -1109 -88 -109
rect 88 -1109 188 -109
rect 364 -1109 464 -109
<< mvndiff >>
rect -522 1097 -464 1109
rect -522 121 -510 1097
rect -476 121 -464 1097
rect -522 109 -464 121
rect -364 1097 -306 1109
rect -364 121 -352 1097
rect -318 121 -306 1097
rect -364 109 -306 121
rect -246 1097 -188 1109
rect -246 121 -234 1097
rect -200 121 -188 1097
rect -246 109 -188 121
rect -88 1097 -30 1109
rect -88 121 -76 1097
rect -42 121 -30 1097
rect -88 109 -30 121
rect 30 1097 88 1109
rect 30 121 42 1097
rect 76 121 88 1097
rect 30 109 88 121
rect 188 1097 246 1109
rect 188 121 200 1097
rect 234 121 246 1097
rect 188 109 246 121
rect 306 1097 364 1109
rect 306 121 318 1097
rect 352 121 364 1097
rect 306 109 364 121
rect 464 1097 522 1109
rect 464 121 476 1097
rect 510 121 522 1097
rect 464 109 522 121
rect -522 -121 -464 -109
rect -522 -1097 -510 -121
rect -476 -1097 -464 -121
rect -522 -1109 -464 -1097
rect -364 -121 -306 -109
rect -364 -1097 -352 -121
rect -318 -1097 -306 -121
rect -364 -1109 -306 -1097
rect -246 -121 -188 -109
rect -246 -1097 -234 -121
rect -200 -1097 -188 -121
rect -246 -1109 -188 -1097
rect -88 -121 -30 -109
rect -88 -1097 -76 -121
rect -42 -1097 -30 -121
rect -88 -1109 -30 -1097
rect 30 -121 88 -109
rect 30 -1097 42 -121
rect 76 -1097 88 -121
rect 30 -1109 88 -1097
rect 188 -121 246 -109
rect 188 -1097 200 -121
rect 234 -1097 246 -121
rect 188 -1109 246 -1097
rect 306 -121 364 -109
rect 306 -1097 318 -121
rect 352 -1097 364 -121
rect 306 -1109 364 -1097
rect 464 -121 522 -109
rect 464 -1097 476 -121
rect 510 -1097 522 -121
rect 464 -1109 522 -1097
<< mvndiffc >>
rect -510 121 -476 1097
rect -352 121 -318 1097
rect -234 121 -200 1097
rect -76 121 -42 1097
rect 42 121 76 1097
rect 200 121 234 1097
rect 318 121 352 1097
rect 476 121 510 1097
rect -510 -1097 -476 -121
rect -352 -1097 -318 -121
rect -234 -1097 -200 -121
rect -76 -1097 -42 -121
rect 42 -1097 76 -121
rect 200 -1097 234 -121
rect 318 -1097 352 -121
rect 476 -1097 510 -121
<< mvpsubdiff >>
rect -656 1319 656 1331
rect -656 1285 -548 1319
rect 548 1285 656 1319
rect -656 1273 656 1285
rect -656 1223 -598 1273
rect -656 -1223 -644 1223
rect -610 -1223 -598 1223
rect 598 1223 656 1273
rect -656 -1273 -598 -1223
rect 598 -1223 610 1223
rect 644 -1223 656 1223
rect 598 -1273 656 -1223
rect -656 -1285 656 -1273
rect -656 -1319 -548 -1285
rect 548 -1319 656 -1285
rect -656 -1331 656 -1319
<< mvpsubdiffcont >>
rect -548 1285 548 1319
rect -644 -1223 -610 1223
rect 610 -1223 644 1223
rect -548 -1319 548 -1285
<< poly >>
rect -464 1181 -364 1197
rect -464 1147 -448 1181
rect -380 1147 -364 1181
rect -464 1109 -364 1147
rect -188 1181 -88 1197
rect -188 1147 -172 1181
rect -104 1147 -88 1181
rect -188 1109 -88 1147
rect 88 1181 188 1197
rect 88 1147 104 1181
rect 172 1147 188 1181
rect 88 1109 188 1147
rect 364 1181 464 1197
rect 364 1147 380 1181
rect 448 1147 464 1181
rect 364 1109 464 1147
rect -464 71 -364 109
rect -464 37 -448 71
rect -380 37 -364 71
rect -464 21 -364 37
rect -188 71 -88 109
rect -188 37 -172 71
rect -104 37 -88 71
rect -188 21 -88 37
rect 88 71 188 109
rect 88 37 104 71
rect 172 37 188 71
rect 88 21 188 37
rect 364 71 464 109
rect 364 37 380 71
rect 448 37 464 71
rect 364 21 464 37
rect -464 -37 -364 -21
rect -464 -71 -448 -37
rect -380 -71 -364 -37
rect -464 -109 -364 -71
rect -188 -37 -88 -21
rect -188 -71 -172 -37
rect -104 -71 -88 -37
rect -188 -109 -88 -71
rect 88 -37 188 -21
rect 88 -71 104 -37
rect 172 -71 188 -37
rect 88 -109 188 -71
rect 364 -37 464 -21
rect 364 -71 380 -37
rect 448 -71 464 -37
rect 364 -109 464 -71
rect -464 -1147 -364 -1109
rect -464 -1181 -448 -1147
rect -380 -1181 -364 -1147
rect -464 -1197 -364 -1181
rect -188 -1147 -88 -1109
rect -188 -1181 -172 -1147
rect -104 -1181 -88 -1147
rect -188 -1197 -88 -1181
rect 88 -1147 188 -1109
rect 88 -1181 104 -1147
rect 172 -1181 188 -1147
rect 88 -1197 188 -1181
rect 364 -1147 464 -1109
rect 364 -1181 380 -1147
rect 448 -1181 464 -1147
rect 364 -1197 464 -1181
<< polycont >>
rect -448 1147 -380 1181
rect -172 1147 -104 1181
rect 104 1147 172 1181
rect 380 1147 448 1181
rect -448 37 -380 71
rect -172 37 -104 71
rect 104 37 172 71
rect 380 37 448 71
rect -448 -71 -380 -37
rect -172 -71 -104 -37
rect 104 -71 172 -37
rect 380 -71 448 -37
rect -448 -1181 -380 -1147
rect -172 -1181 -104 -1147
rect 104 -1181 172 -1147
rect 380 -1181 448 -1147
<< locali >>
rect -644 1285 -548 1319
rect 548 1285 644 1319
rect -644 1223 -610 1285
rect 610 1223 644 1285
rect -464 1147 -448 1181
rect -380 1147 -364 1181
rect -188 1147 -172 1181
rect -104 1147 -88 1181
rect 88 1147 104 1181
rect 172 1147 188 1181
rect 364 1147 380 1181
rect 448 1147 464 1181
rect -510 1097 -476 1113
rect -510 105 -476 121
rect -352 1097 -318 1113
rect -352 105 -318 121
rect -234 1097 -200 1113
rect -234 105 -200 121
rect -76 1097 -42 1113
rect -76 105 -42 121
rect 42 1097 76 1113
rect 42 105 76 121
rect 200 1097 234 1113
rect 200 105 234 121
rect 318 1097 352 1113
rect 318 105 352 121
rect 476 1097 510 1113
rect 476 105 510 121
rect -464 37 -448 71
rect -380 37 -364 71
rect -188 37 -172 71
rect -104 37 -88 71
rect 88 37 104 71
rect 172 37 188 71
rect 364 37 380 71
rect 448 37 464 71
rect -464 -71 -448 -37
rect -380 -71 -364 -37
rect -188 -71 -172 -37
rect -104 -71 -88 -37
rect 88 -71 104 -37
rect 172 -71 188 -37
rect 364 -71 380 -37
rect 448 -71 464 -37
rect -510 -121 -476 -105
rect -510 -1113 -476 -1097
rect -352 -121 -318 -105
rect -352 -1113 -318 -1097
rect -234 -121 -200 -105
rect -234 -1113 -200 -1097
rect -76 -121 -42 -105
rect -76 -1113 -42 -1097
rect 42 -121 76 -105
rect 42 -1113 76 -1097
rect 200 -121 234 -105
rect 200 -1113 234 -1097
rect 318 -121 352 -105
rect 318 -1113 352 -1097
rect 476 -121 510 -105
rect 476 -1113 510 -1097
rect -464 -1181 -448 -1147
rect -380 -1181 -364 -1147
rect -188 -1181 -172 -1147
rect -104 -1181 -88 -1147
rect 88 -1181 104 -1147
rect 172 -1181 188 -1147
rect 364 -1181 380 -1147
rect 448 -1181 464 -1147
rect -644 -1285 -610 -1223
rect 610 -1285 644 -1223
rect -644 -1319 -548 -1285
rect 548 -1319 644 -1285
<< viali >>
rect -448 1147 -380 1181
rect -172 1147 -104 1181
rect 104 1147 172 1181
rect 380 1147 448 1181
rect -510 121 -476 1097
rect -352 121 -318 1097
rect -234 121 -200 1097
rect -76 121 -42 1097
rect 42 121 76 1097
rect 200 121 234 1097
rect 318 121 352 1097
rect 476 121 510 1097
rect -448 37 -380 71
rect -172 37 -104 71
rect 104 37 172 71
rect 380 37 448 71
rect -448 -71 -380 -37
rect -172 -71 -104 -37
rect 104 -71 172 -37
rect 380 -71 448 -37
rect -510 -1097 -476 -121
rect -352 -1097 -318 -121
rect -234 -1097 -200 -121
rect -76 -1097 -42 -121
rect 42 -1097 76 -121
rect 200 -1097 234 -121
rect 318 -1097 352 -121
rect 476 -1097 510 -121
rect -448 -1181 -380 -1147
rect -172 -1181 -104 -1147
rect 104 -1181 172 -1147
rect 380 -1181 448 -1147
<< metal1 >>
rect -460 1181 -368 1187
rect -460 1147 -448 1181
rect -380 1147 -368 1181
rect -460 1141 -368 1147
rect -184 1181 -92 1187
rect -184 1147 -172 1181
rect -104 1147 -92 1181
rect -184 1141 -92 1147
rect 92 1181 184 1187
rect 92 1147 104 1181
rect 172 1147 184 1181
rect 92 1141 184 1147
rect 368 1181 460 1187
rect 368 1147 380 1181
rect 448 1147 460 1181
rect 368 1141 460 1147
rect -516 1097 -470 1109
rect -516 121 -510 1097
rect -476 121 -470 1097
rect -516 109 -470 121
rect -358 1097 -312 1109
rect -358 121 -352 1097
rect -318 121 -312 1097
rect -358 109 -312 121
rect -240 1097 -194 1109
rect -240 121 -234 1097
rect -200 121 -194 1097
rect -240 109 -194 121
rect -82 1097 -36 1109
rect -82 121 -76 1097
rect -42 121 -36 1097
rect -82 109 -36 121
rect 36 1097 82 1109
rect 36 121 42 1097
rect 76 121 82 1097
rect 36 109 82 121
rect 194 1097 240 1109
rect 194 121 200 1097
rect 234 121 240 1097
rect 194 109 240 121
rect 312 1097 358 1109
rect 312 121 318 1097
rect 352 121 358 1097
rect 312 109 358 121
rect 470 1097 516 1109
rect 470 121 476 1097
rect 510 121 516 1097
rect 470 109 516 121
rect -460 71 -368 77
rect -460 37 -448 71
rect -380 37 -368 71
rect -460 31 -368 37
rect -184 71 -92 77
rect -184 37 -172 71
rect -104 37 -92 71
rect -184 31 -92 37
rect 92 71 184 77
rect 92 37 104 71
rect 172 37 184 71
rect 92 31 184 37
rect 368 71 460 77
rect 368 37 380 71
rect 448 37 460 71
rect 368 31 460 37
rect -460 -37 -368 -31
rect -460 -71 -448 -37
rect -380 -71 -368 -37
rect -460 -77 -368 -71
rect -184 -37 -92 -31
rect -184 -71 -172 -37
rect -104 -71 -92 -37
rect -184 -77 -92 -71
rect 92 -37 184 -31
rect 92 -71 104 -37
rect 172 -71 184 -37
rect 92 -77 184 -71
rect 368 -37 460 -31
rect 368 -71 380 -37
rect 448 -71 460 -37
rect 368 -77 460 -71
rect -516 -121 -470 -109
rect -516 -1097 -510 -121
rect -476 -1097 -470 -121
rect -516 -1109 -470 -1097
rect -358 -121 -312 -109
rect -358 -1097 -352 -121
rect -318 -1097 -312 -121
rect -358 -1109 -312 -1097
rect -240 -121 -194 -109
rect -240 -1097 -234 -121
rect -200 -1097 -194 -121
rect -240 -1109 -194 -1097
rect -82 -121 -36 -109
rect -82 -1097 -76 -121
rect -42 -1097 -36 -121
rect -82 -1109 -36 -1097
rect 36 -121 82 -109
rect 36 -1097 42 -121
rect 76 -1097 82 -121
rect 36 -1109 82 -1097
rect 194 -121 240 -109
rect 194 -1097 200 -121
rect 234 -1097 240 -121
rect 194 -1109 240 -1097
rect 312 -121 358 -109
rect 312 -1097 318 -121
rect 352 -1097 358 -121
rect 312 -1109 358 -1097
rect 470 -121 516 -109
rect 470 -1097 476 -121
rect 510 -1097 516 -121
rect 470 -1109 516 -1097
rect -460 -1147 -368 -1141
rect -460 -1181 -448 -1147
rect -380 -1181 -368 -1147
rect -460 -1187 -368 -1181
rect -184 -1147 -92 -1141
rect -184 -1181 -172 -1147
rect -104 -1181 -92 -1147
rect -184 -1187 -92 -1181
rect 92 -1147 184 -1141
rect 92 -1181 104 -1147
rect 172 -1181 184 -1147
rect 92 -1187 184 -1181
rect 368 -1147 460 -1141
rect 368 -1181 380 -1147
rect 448 -1181 460 -1147
rect 368 -1187 460 -1181
<< properties >>
string gencell sky130_fd_pr__nfet_03v3_nvt
string FIXED_BBOX -627 -1302 627 1302
string parameters w 5 l 0.50 m 2 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
