magic
tech sky130A
magscale 1 2
timestamp 1697652271
<< pwell >>
rect -201 -1018 201 1018
<< psubdiff >>
rect -165 948 -69 982
rect 69 948 165 982
rect -165 886 -131 948
rect 131 886 165 948
rect -165 -948 -131 -886
rect 131 -948 165 -886
rect -165 -982 -69 -948
rect 69 -982 165 -948
<< psubdiffcont >>
rect -69 948 69 982
rect -165 -886 -131 886
rect 131 -886 165 886
rect -69 -982 69 -948
<< xpolycontact >>
rect -35 420 35 852
rect -35 -852 35 -420
<< xpolyres >>
rect -35 -420 35 420
<< locali >>
rect -165 948 -69 982
rect 69 948 165 982
rect -165 886 -131 948
rect 131 886 165 948
rect -165 -948 -131 -886
rect 131 -948 165 -886
rect -165 -982 -69 -948
rect 69 -982 165 -948
<< viali >>
rect -19 437 19 834
rect -19 -834 19 -437
<< metal1 >>
rect -25 834 25 846
rect -25 437 -19 834
rect 19 437 25 834
rect -25 425 25 437
rect -25 -437 25 -425
rect -25 -834 -19 -437
rect 19 -834 25 -437
rect -25 -846 25 -834
<< res0p35 >>
rect -37 -422 37 422
<< properties >>
string FIXED_BBOX -148 -965 148 965
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 4.2 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 25.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
