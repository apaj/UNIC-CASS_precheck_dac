magic
tech sky130A
magscale 1 2
timestamp 1698012353
<< pwell >>
rect -235 -1228 235 1228
<< psubdiff >>
rect -199 1158 -103 1192
rect 103 1158 199 1192
rect -199 1096 -165 1158
rect 165 1096 199 1158
rect -199 -1158 -165 -1096
rect 165 -1158 199 -1096
rect -199 -1192 -103 -1158
rect 103 -1192 199 -1158
<< psubdiffcont >>
rect -103 1158 103 1192
rect -199 -1096 -165 1096
rect 165 -1096 199 1096
rect -103 -1192 103 -1158
<< xpolycontact >>
rect -69 630 69 1062
rect -69 -1062 69 -630
<< xpolyres >>
rect -69 -630 69 630
<< locali >>
rect -199 1158 -103 1192
rect 103 1158 199 1192
rect -199 1096 -165 1158
rect 165 1096 199 1158
rect -199 -1158 -165 -1096
rect 165 -1158 199 -1096
rect -199 -1192 -103 -1158
rect 103 -1192 199 -1158
<< viali >>
rect -53 647 53 1044
rect -53 -1044 53 -647
<< metal1 >>
rect -59 1044 59 1056
rect -59 647 -53 1044
rect 53 647 59 1044
rect -59 635 59 647
rect -59 -647 59 -635
rect -59 -1044 -53 -647
rect 53 -1044 59 -647
rect -59 -1056 59 -1044
<< res0p69 >>
rect -71 -632 71 632
<< properties >>
string FIXED_BBOX -182 -1175 182 1175
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 6.3 m 1 nx 1 wmin 0.690 lmin 0.50 rho 2000 val 18.806k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
