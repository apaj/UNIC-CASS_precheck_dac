magic
tech sky130A
magscale 1 2
timestamp 1628499526
<< pwell >>
rect -278 -5603 278 5603
<< mvnmos >>
rect -50 3745 50 5345
rect -50 1927 50 3527
rect -50 109 50 1709
rect -50 -1709 50 -109
rect -50 -3527 50 -1927
rect -50 -5345 50 -3745
<< mvndiff >>
rect -108 5333 -50 5345
rect -108 3757 -96 5333
rect -62 3757 -50 5333
rect -108 3745 -50 3757
rect 50 5333 108 5345
rect 50 3757 62 5333
rect 96 3757 108 5333
rect 50 3745 108 3757
rect -108 3515 -50 3527
rect -108 1939 -96 3515
rect -62 1939 -50 3515
rect -108 1927 -50 1939
rect 50 3515 108 3527
rect 50 1939 62 3515
rect 96 1939 108 3515
rect 50 1927 108 1939
rect -108 1697 -50 1709
rect -108 121 -96 1697
rect -62 121 -50 1697
rect -108 109 -50 121
rect 50 1697 108 1709
rect 50 121 62 1697
rect 96 121 108 1697
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -1697 -96 -121
rect -62 -1697 -50 -121
rect -108 -1709 -50 -1697
rect 50 -121 108 -109
rect 50 -1697 62 -121
rect 96 -1697 108 -121
rect 50 -1709 108 -1697
rect -108 -1939 -50 -1927
rect -108 -3515 -96 -1939
rect -62 -3515 -50 -1939
rect -108 -3527 -50 -3515
rect 50 -1939 108 -1927
rect 50 -3515 62 -1939
rect 96 -3515 108 -1939
rect 50 -3527 108 -3515
rect -108 -3757 -50 -3745
rect -108 -5333 -96 -3757
rect -62 -5333 -50 -3757
rect -108 -5345 -50 -5333
rect 50 -3757 108 -3745
rect 50 -5333 62 -3757
rect 96 -5333 108 -3757
rect 50 -5345 108 -5333
<< mvndiffc >>
rect -96 3757 -62 5333
rect 62 3757 96 5333
rect -96 1939 -62 3515
rect 62 1939 96 3515
rect -96 121 -62 1697
rect 62 121 96 1697
rect -96 -1697 -62 -121
rect 62 -1697 96 -121
rect -96 -3515 -62 -1939
rect 62 -3515 96 -1939
rect -96 -5333 -62 -3757
rect 62 -5333 96 -3757
<< mvpsubdiff >>
rect -242 5555 242 5567
rect -242 5521 -134 5555
rect 134 5521 242 5555
rect -242 5509 242 5521
rect -242 5459 -184 5509
rect -242 -5459 -230 5459
rect -196 -5459 -184 5459
rect 184 5459 242 5509
rect -242 -5509 -184 -5459
rect 184 -5459 196 5459
rect 230 -5459 242 5459
rect 184 -5509 242 -5459
rect -242 -5521 242 -5509
rect -242 -5555 -134 -5521
rect 134 -5555 242 -5521
rect -242 -5567 242 -5555
<< mvpsubdiffcont >>
rect -134 5521 134 5555
rect -230 -5459 -196 5459
rect 196 -5459 230 5459
rect -134 -5555 134 -5521
<< poly >>
rect -50 5417 50 5433
rect -50 5383 -34 5417
rect 34 5383 50 5417
rect -50 5345 50 5383
rect -50 3707 50 3745
rect -50 3673 -34 3707
rect 34 3673 50 3707
rect -50 3657 50 3673
rect -50 3599 50 3615
rect -50 3565 -34 3599
rect 34 3565 50 3599
rect -50 3527 50 3565
rect -50 1889 50 1927
rect -50 1855 -34 1889
rect 34 1855 50 1889
rect -50 1839 50 1855
rect -50 1781 50 1797
rect -50 1747 -34 1781
rect 34 1747 50 1781
rect -50 1709 50 1747
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -1747 50 -1709
rect -50 -1781 -34 -1747
rect 34 -1781 50 -1747
rect -50 -1797 50 -1781
rect -50 -1855 50 -1839
rect -50 -1889 -34 -1855
rect 34 -1889 50 -1855
rect -50 -1927 50 -1889
rect -50 -3565 50 -3527
rect -50 -3599 -34 -3565
rect 34 -3599 50 -3565
rect -50 -3615 50 -3599
rect -50 -3673 50 -3657
rect -50 -3707 -34 -3673
rect 34 -3707 50 -3673
rect -50 -3745 50 -3707
rect -50 -5383 50 -5345
rect -50 -5417 -34 -5383
rect 34 -5417 50 -5383
rect -50 -5433 50 -5417
<< polycont >>
rect -34 5383 34 5417
rect -34 3673 34 3707
rect -34 3565 34 3599
rect -34 1855 34 1889
rect -34 1747 34 1781
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -1781 34 -1747
rect -34 -1889 34 -1855
rect -34 -3599 34 -3565
rect -34 -3707 34 -3673
rect -34 -5417 34 -5383
<< locali >>
rect -230 5521 -134 5555
rect 134 5521 230 5555
rect -230 5459 -196 5521
rect 196 5459 230 5521
rect -50 5383 -34 5417
rect 34 5383 50 5417
rect -96 5333 -62 5349
rect -96 3741 -62 3757
rect 62 5333 96 5349
rect 62 3741 96 3757
rect -50 3673 -34 3707
rect 34 3673 50 3707
rect -50 3565 -34 3599
rect 34 3565 50 3599
rect -96 3515 -62 3531
rect -96 1923 -62 1939
rect 62 3515 96 3531
rect 62 1923 96 1939
rect -50 1855 -34 1889
rect 34 1855 50 1889
rect -50 1747 -34 1781
rect 34 1747 50 1781
rect -96 1697 -62 1713
rect -96 105 -62 121
rect 62 1697 96 1713
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -1713 -62 -1697
rect 62 -121 96 -105
rect 62 -1713 96 -1697
rect -50 -1781 -34 -1747
rect 34 -1781 50 -1747
rect -50 -1889 -34 -1855
rect 34 -1889 50 -1855
rect -96 -1939 -62 -1923
rect -96 -3531 -62 -3515
rect 62 -1939 96 -1923
rect 62 -3531 96 -3515
rect -50 -3599 -34 -3565
rect 34 -3599 50 -3565
rect -50 -3707 -34 -3673
rect 34 -3707 50 -3673
rect -96 -3757 -62 -3741
rect -96 -5349 -62 -5333
rect 62 -3757 96 -3741
rect 62 -5349 96 -5333
rect -50 -5417 -34 -5383
rect 34 -5417 50 -5383
rect -230 -5521 -196 -5459
rect 196 -5521 230 -5459
rect -230 -5555 -134 -5521
rect 134 -5555 230 -5521
<< viali >>
rect -34 5383 34 5417
rect -96 3757 -62 5333
rect 62 3757 96 5333
rect -34 3673 34 3707
rect -34 3565 34 3599
rect -96 1939 -62 3515
rect 62 1939 96 3515
rect -34 1855 34 1889
rect -34 1747 34 1781
rect -96 121 -62 1697
rect 62 121 96 1697
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -1697 -62 -121
rect 62 -1697 96 -121
rect -34 -1781 34 -1747
rect -34 -1889 34 -1855
rect -96 -3515 -62 -1939
rect 62 -3515 96 -1939
rect -34 -3599 34 -3565
rect -34 -3707 34 -3673
rect -96 -5333 -62 -3757
rect 62 -5333 96 -3757
rect -34 -5417 34 -5383
<< metal1 >>
rect -46 5417 46 5423
rect -46 5383 -34 5417
rect 34 5383 46 5417
rect -46 5377 46 5383
rect -102 5333 -56 5345
rect -102 3757 -96 5333
rect -62 3757 -56 5333
rect -102 3745 -56 3757
rect 56 5333 102 5345
rect 56 3757 62 5333
rect 96 3757 102 5333
rect 56 3745 102 3757
rect -46 3707 46 3713
rect -46 3673 -34 3707
rect 34 3673 46 3707
rect -46 3667 46 3673
rect -46 3599 46 3605
rect -46 3565 -34 3599
rect 34 3565 46 3599
rect -46 3559 46 3565
rect -102 3515 -56 3527
rect -102 1939 -96 3515
rect -62 1939 -56 3515
rect -102 1927 -56 1939
rect 56 3515 102 3527
rect 56 1939 62 3515
rect 96 1939 102 3515
rect 56 1927 102 1939
rect -46 1889 46 1895
rect -46 1855 -34 1889
rect 34 1855 46 1889
rect -46 1849 46 1855
rect -46 1781 46 1787
rect -46 1747 -34 1781
rect 34 1747 46 1781
rect -46 1741 46 1747
rect -102 1697 -56 1709
rect -102 121 -96 1697
rect -62 121 -56 1697
rect -102 109 -56 121
rect 56 1697 102 1709
rect 56 121 62 1697
rect 96 121 102 1697
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -1697 -96 -121
rect -62 -1697 -56 -121
rect -102 -1709 -56 -1697
rect 56 -121 102 -109
rect 56 -1697 62 -121
rect 96 -1697 102 -121
rect 56 -1709 102 -1697
rect -46 -1747 46 -1741
rect -46 -1781 -34 -1747
rect 34 -1781 46 -1747
rect -46 -1787 46 -1781
rect -46 -1855 46 -1849
rect -46 -1889 -34 -1855
rect 34 -1889 46 -1855
rect -46 -1895 46 -1889
rect -102 -1939 -56 -1927
rect -102 -3515 -96 -1939
rect -62 -3515 -56 -1939
rect -102 -3527 -56 -3515
rect 56 -1939 102 -1927
rect 56 -3515 62 -1939
rect 96 -3515 102 -1939
rect 56 -3527 102 -3515
rect -46 -3565 46 -3559
rect -46 -3599 -34 -3565
rect 34 -3599 46 -3565
rect -46 -3605 46 -3599
rect -46 -3673 46 -3667
rect -46 -3707 -34 -3673
rect 34 -3707 46 -3673
rect -46 -3713 46 -3707
rect -102 -3757 -56 -3745
rect -102 -5333 -96 -3757
rect -62 -5333 -56 -3757
rect -102 -5345 -56 -5333
rect 56 -3757 102 -3745
rect 56 -5333 62 -3757
rect 96 -5333 102 -3757
rect 56 -5345 102 -5333
rect -46 -5383 46 -5377
rect -46 -5417 -34 -5383
rect 34 -5417 46 -5383
rect -46 -5423 46 -5417
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -213 -5538 213 5538
string parameters w 8 l 0.50 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
