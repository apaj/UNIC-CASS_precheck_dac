* SPICE3 file created from dac_cell2.ext - technology: sky130A

.option scale=5000u

.subckt dac_cell2 vsup vgnd iref vsw iout iout_n vbias
X0 m1_4330_3580# m1_n2460_3700# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=5400
X1 m1_4330_3580# m1_n2460_3700# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=5400
X2 m1_4330_3580# vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=5400
X3 m1_4330_3580# vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=5400
X4 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 ad=11600 pd=516 as=11600 ps=516 w=200 l=200
X5 m1_n1250_930# iref m1_n2460_3700# vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=400 l=200
X6 iout vsw m1_n1250_930# vsup sky130_fd_pr__pfet_g5v0d10v5 ad=23200 pd=916 as=0 ps=0 w=400 l=200
X7 iout_n vbias m1_n1250_930# vsup sky130_fd_pr__pfet_g5v0d10v5 ad=23200 pd=916 as=0 ps=0 w=400 l=200
.ends
