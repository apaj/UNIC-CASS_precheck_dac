magic
tech sky130A
magscale 1 2
timestamp 1698012353
<< viali >>
rect 4860 5000 4900 5210
rect 4860 4510 4910 4720
rect 4860 4020 4900 4230
rect 4850 3540 4890 3750
rect -1810 2220 -1450 2260
rect -690 2130 -310 2180
rect -700 1520 -320 1560
rect 480 1520 860 1560
<< metal1 >>
rect 4800 5210 5000 5250
rect -1510 5000 -1070 5180
rect -2930 4930 -1070 5000
rect -3290 4740 -1070 4930
rect -3290 4730 -2570 4740
rect -2920 2640 -2570 4730
rect -1510 4560 -1070 4740
rect -1490 4060 -1050 4190
rect -2460 4010 -1050 4060
rect -2460 3780 -2400 4010
rect -2160 3780 -1050 4010
rect -2460 3700 -1050 3780
rect -1490 3570 -1050 3700
rect 4330 3580 4770 5180
rect 4800 5000 4860 5210
rect 4900 5000 5000 5210
rect 4800 4720 5000 5000
rect 4800 4510 4860 4720
rect 4910 4510 5000 4720
rect 4800 4230 5000 4510
rect 4800 4020 4860 4230
rect 4900 4020 5000 4230
rect 4800 3750 5000 4020
rect 4800 3540 4850 3750
rect 4890 3540 5000 3750
rect 4800 3140 5000 3540
rect -1730 2800 -410 2910
rect -1730 2680 -1540 2800
rect -2920 2430 -1740 2640
rect -1130 2630 -990 2800
rect -1520 2610 -990 2630
rect -1520 2480 -1380 2610
rect -1210 2480 -990 2610
rect -1520 2450 -990 2480
rect -900 2680 -620 2750
rect -900 2450 -860 2680
rect -690 2450 -620 2680
rect -2920 2420 -2430 2430
rect -2580 2210 -2430 2420
rect -900 2360 -620 2450
rect -390 2680 290 2720
rect -390 2410 -30 2680
rect 240 2410 290 2680
rect 4800 2550 5010 3140
rect -390 2380 290 2410
rect -1830 2260 -1430 2280
rect -1830 2220 -1810 2260
rect -1450 2220 -1430 2260
rect -1830 2210 -1430 2220
rect -2580 2180 -290 2210
rect -2580 2130 -690 2180
rect -310 2130 -290 2180
rect -2580 2110 -290 2130
rect -2520 1890 -2320 1900
rect -2520 1510 -2320 1760
rect -720 1590 -290 2110
rect -720 1560 870 1590
rect -720 1520 -700 1560
rect -320 1520 480 1560
rect 860 1520 870 1560
rect -720 1500 870 1520
rect -1250 1240 -620 1330
rect -1250 1000 -1200 1240
rect -970 1000 -620 1240
rect -1250 950 -620 1000
rect -400 950 -120 1330
rect -1250 930 -630 950
rect -610 410 -420 890
rect -280 520 -120 950
rect -40 1260 560 1330
rect -40 1020 40 1260
rect 290 1020 560 1260
rect -40 940 560 1020
rect 780 950 1310 1330
rect -610 70 -410 410
rect -280 320 210 520
rect 570 440 760 900
rect 1100 550 1310 950
rect 570 40 770 440
rect 1100 350 1800 550
<< via1 >>
rect -2400 3780 -2160 4010
rect -1380 2480 -1210 2610
rect -860 2450 -690 2680
rect -30 2410 240 2680
rect -2520 1760 -2320 1890
rect -1200 1000 -970 1240
rect 40 1020 290 1260
<< metal2 >>
rect -2470 4010 -2140 4030
rect -2470 3780 -2400 4010
rect -2160 3780 -2140 4010
rect -2470 3220 -2140 3780
rect -2470 3020 -880 3220
rect -1150 2710 -880 3020
rect -1150 2680 -660 2710
rect -1420 2610 -1180 2650
rect -1420 2480 -1380 2610
rect -1210 2480 -1180 2610
rect -1420 2060 -1180 2480
rect -1150 2450 -860 2680
rect -690 2450 -660 2680
rect -1150 2440 -660 2450
rect -890 2420 -660 2440
rect -100 2680 300 2720
rect -2540 1920 -1180 2060
rect -100 2410 -30 2680
rect 240 2410 300 2680
rect -2540 1890 -2280 1920
rect -2540 1760 -2520 1890
rect -2320 1760 -2280 1890
rect -100 1870 300 2410
rect -2540 1740 -2280 1760
rect -1250 1690 300 1870
rect -1250 1330 -960 1690
rect -1250 1240 -930 1330
rect 10 1300 300 1690
rect -1250 1000 -1200 1240
rect -970 1000 -930 1240
rect -1250 930 -930 1000
rect -30 1260 320 1300
rect -30 1020 40 1260
rect 290 1020 320 1260
rect -30 950 320 1020
use sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#1  XM1
timestamp 1698012353
transform 1 0 -1632 0 1 2537
box -358 -397 358 397
use sky130_fd_pr__pfet_g5v0d10v5_FGK6VM  XM2
timestamp 1698012353
transform 1 0 -502 0 1 2557
box -358 -497 358 497
use sky130_fd_pr__pfet_g5v0d10v5_FGK6VM  XM3
timestamp 1698012353
transform 1 0 -512 0 1 1137
box -358 -497 358 497
use sky130_fd_pr__pfet_g5v0d10v5_FGK6VM  XM4
timestamp 1698012353
transform 1 0 668 0 1 1137
box -358 -497 358 497
use sky130_fd_pr__res_xhigh_po_0p69_XZX24Q  XR1
timestamp 1698012353
transform 0 -1 1628 1 0 3645
box -235 -3298 235 3298
use sky130_fd_pr__res_xhigh_po_0p69_XZX24Q  XR2
timestamp 1698012353
transform 0 -1 1638 1 0 4125
box -235 -3298 235 3298
use sky130_fd_pr__res_xhigh_po_0p69_XZX24Q  XR3
timestamp 1698012353
transform 0 -1 1638 1 0 4615
box -235 -3298 235 3298
use sky130_fd_pr__res_xhigh_po_0p69_XZX24Q  XR4
timestamp 1698012353
transform 0 -1 1638 1 0 5105
box -235 -3298 235 3298
<< labels >>
flabel metal1 -3290 4730 -3090 4930 0 FreeSans 1280 0 0 0 vsup
port 0 nsew
flabel metal1 4810 2550 5010 2750 0 FreeSans 1280 0 0 0 vgnd
port 1 nsew
flabel metal1 10 320 210 520 0 FreeSans 1280 0 0 0 iout
port 4 nsew
flabel metal1 1600 350 1800 550 0 FreeSans 1280 0 0 0 iout_n
port 5 nsew
flabel metal1 -610 70 -410 270 0 FreeSans 1280 0 0 0 vsw
port 3 nsew
flabel metal1 570 40 770 240 0 FreeSans 1280 0 0 0 vbias
port 6 nsew
flabel metal1 -2520 1510 -2320 1710 0 FreeSans 1280 0 0 0 iref
port 2 nsew
rlabel metal2 -92 1816 276 1996 1 sourceM3M4
rlabel metal2 -1576 3032 -1208 3212 1 sourceM2
rlabel metal1 4396 4020 4648 4660 1 parR
<< end >>
