* NGSPICE file created from dac_cell2.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p69_XZX24Q a_n199_n3262# a_n69_n3132# a_n69_2700#
X0 a_n69_2700# a_n69_n3132# a_n199_n3262# sky130_fd_pr__res_xhigh_po_0p69 l=27
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#1 a_n100_n197# a_100_n100# w_n358_n397#
+ a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n358_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGK6VM a_n100_n297# a_100_n200# w_n358_n497#
+ a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n358_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt dac_cell2 vsup vgnd iref vsw iout iout_n vbias
XXR1 vgnd parR sourceM2 sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR2 vgnd parR sourceM2 sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR3 vgnd parR vsup sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR4 vgnd parR vsup sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#1
XXM2 iref sourceM3M4 vsup sourceM2 sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
XXM3 vsw iout vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
XXM4 vbias iout_n vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
.ends

