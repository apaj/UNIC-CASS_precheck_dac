magic
tech sky130A
magscale 1 2
timestamp 1697533315
<< nwell >>
rect -466 -997 466 997
<< mvpmos >>
rect -208 -700 -108 700
rect -50 -700 50 700
rect 108 -700 208 700
<< mvpdiff >>
rect -266 688 -208 700
rect -266 -688 -254 688
rect -220 -688 -208 688
rect -266 -700 -208 -688
rect -108 688 -50 700
rect -108 -688 -96 688
rect -62 -688 -50 688
rect -108 -700 -50 -688
rect 50 688 108 700
rect 50 -688 62 688
rect 96 -688 108 688
rect 50 -700 108 -688
rect 208 688 266 700
rect 208 -688 220 688
rect 254 -688 266 688
rect 208 -700 266 -688
<< mvpdiffc >>
rect -254 -688 -220 688
rect -96 -688 -62 688
rect 62 -688 96 688
rect 220 -688 254 688
<< mvnsubdiff >>
rect -400 919 400 931
rect -400 885 -292 919
rect 292 885 400 919
rect -400 873 400 885
rect -400 823 -342 873
rect -400 -823 -388 823
rect -354 -823 -342 823
rect 342 823 400 873
rect -400 -873 -342 -823
rect 342 -823 354 823
rect 388 -823 400 823
rect 342 -873 400 -823
rect -400 -885 400 -873
rect -400 -919 -292 -885
rect 292 -919 400 -885
rect -400 -931 400 -919
<< mvnsubdiffcont >>
rect -292 885 292 919
rect -388 -823 -354 823
rect 354 -823 388 823
rect -292 -919 292 -885
<< poly >>
rect -208 781 -108 797
rect -208 747 -192 781
rect -124 747 -108 781
rect -208 700 -108 747
rect -50 781 50 797
rect -50 747 -34 781
rect 34 747 50 781
rect -50 700 50 747
rect 108 781 208 797
rect 108 747 124 781
rect 192 747 208 781
rect 108 700 208 747
rect -208 -747 -108 -700
rect -208 -781 -192 -747
rect -124 -781 -108 -747
rect -208 -797 -108 -781
rect -50 -747 50 -700
rect -50 -781 -34 -747
rect 34 -781 50 -747
rect -50 -797 50 -781
rect 108 -747 208 -700
rect 108 -781 124 -747
rect 192 -781 208 -747
rect 108 -797 208 -781
<< polycont >>
rect -192 747 -124 781
rect -34 747 34 781
rect 124 747 192 781
rect -192 -781 -124 -747
rect -34 -781 34 -747
rect 124 -781 192 -747
<< locali >>
rect -388 885 -292 919
rect 292 885 388 919
rect -388 823 -354 885
rect 354 823 388 885
rect -208 747 -192 781
rect -124 747 -108 781
rect -50 747 -34 781
rect 34 747 50 781
rect 108 747 124 781
rect 192 747 208 781
rect -254 688 -220 704
rect -254 -704 -220 -688
rect -96 688 -62 704
rect -96 -704 -62 -688
rect 62 688 96 704
rect 62 -704 96 -688
rect 220 688 254 704
rect 220 -704 254 -688
rect -208 -781 -192 -747
rect -124 -781 -108 -747
rect -50 -781 -34 -747
rect 34 -781 50 -747
rect 108 -781 124 -747
rect 192 -781 208 -747
rect -388 -885 -354 -823
rect 354 -885 388 -823
rect -388 -919 -292 -885
rect 292 -919 388 -885
<< viali >>
rect -192 747 -124 781
rect -34 747 34 781
rect 124 747 192 781
rect -254 -688 -220 688
rect -96 -688 -62 688
rect 62 -688 96 688
rect 220 -688 254 688
rect -192 -781 -124 -747
rect -34 -781 34 -747
rect 124 -781 192 -747
<< metal1 >>
rect -204 781 -112 787
rect -204 747 -192 781
rect -124 747 -112 781
rect -204 741 -112 747
rect -46 781 46 787
rect -46 747 -34 781
rect 34 747 46 781
rect -46 741 46 747
rect 112 781 204 787
rect 112 747 124 781
rect 192 747 204 781
rect 112 741 204 747
rect -260 688 -214 700
rect -260 -688 -254 688
rect -220 -688 -214 688
rect -260 -700 -214 -688
rect -102 688 -56 700
rect -102 -688 -96 688
rect -62 -688 -56 688
rect -102 -700 -56 -688
rect 56 688 102 700
rect 56 -688 62 688
rect 96 -688 102 688
rect 56 -700 102 -688
rect 214 688 260 700
rect 214 -688 220 688
rect 254 -688 260 688
rect 214 -700 260 -688
rect -204 -747 -112 -741
rect -204 -781 -192 -747
rect -124 -781 -112 -747
rect -204 -787 -112 -781
rect -46 -747 46 -741
rect -46 -781 -34 -747
rect 34 -781 46 -747
rect -46 -787 46 -781
rect 112 -747 204 -741
rect 112 -781 124 -747
rect 192 -781 204 -747
rect 112 -787 204 -781
<< properties >>
string FIXED_BBOX -371 -902 371 902
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 7.0 l 0.5 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
