**.subckt tb_dac_cell1_tran
V1 net5 GND 3.3
V2 Vsw GND pulse(0, 3.3, 20ms, 1ns, 1ns, 10ms, 20ms)
V3 net6 GND 0.7
V4 net7 net3 0
V5 net2 net1 0
R1 net1 GND 200 m=1
R2 net3 GND 200 m=1
R4 net4 GND 150k m=1
x1 net5 net4 GND Vsw net6 net7 net2 dac_cell1
**** begin user architecture code


.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.param mc_pr_switch=0
*** ANALYSIS TO DO

.tran 0.1 150m 0.001m
.save i(V4) i(V5)
.save Vsw

.control
set wr_vecnames
set wr_singlescale

run
******** results filename  ************ nodes to write
wrdata $DEV_PATH/res/dac_cell1_tran_cur.res i(V4) i(V5)
wrdata $DEV_PATH/res/dac_cell1_tran_vol.res Vsw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  dac_cell1.sym # of pins=7
* sym_path: /opt/uniccass/dev/dac_cell1/tb/dac_cell1.sym
* sch_path: /opt/uniccass/dev/dac_cell1/tb/dac_cell1.sch
.subckt dac_cell1  vsup iref vgnd vsw vbias iout_n iout
*.iopin vsup
*.iopin vgnd
*.iopin iref
*.iopin vsw
*.iopin iout
*.iopin iout_n
*.iopin vbias
XM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 sourceM3M4 iref sourceM2 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 iout vsw sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 iout_n vbias sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XR1 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
XR2 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
XR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
XR4 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
.ends

.GLOBAL GND
** flattened .save nodes
.save i(V4) i(V5)
.save Vsw
.end
