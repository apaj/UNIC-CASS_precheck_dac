magic
tech sky130A
magscale 1 2
timestamp 1695199131
<< viali >>
rect 1132 6906 1180 7272
rect 78 508 528 544
rect 1686 74 1730 442
rect 1708 -938 1744 -566
rect 2152 -958 2188 -586
<< metal1 >>
rect 1170 14168 1622 14414
rect 200 14118 2430 14168
rect 200 13802 2436 14118
rect 200 7278 384 13802
rect 2104 13214 2436 13802
rect 1302 13062 3210 13214
rect 1322 7654 3230 7806
rect 2094 7364 2432 7654
rect 1124 7278 1186 7284
rect 200 7272 1186 7278
rect 200 6906 1132 7272
rect 1180 6906 1186 7272
rect 1312 7212 3220 7364
rect 200 6902 1186 6906
rect 200 2912 384 6902
rect 1124 6894 1186 6902
rect 200 2852 390 2912
rect 204 1704 390 2852
rect 1296 1788 3204 1940
rect 204 1584 392 1704
rect 206 932 392 1584
rect 2100 1364 2438 1788
rect 1312 1342 2438 1364
rect 1312 1288 2436 1342
rect 206 688 214 932
rect 380 688 392 932
rect 206 558 392 688
rect 1310 1132 2436 1288
rect 56 544 548 558
rect 56 508 78 544
rect 528 508 548 544
rect 56 496 548 508
rect 206 376 392 496
rect 434 170 1280 356
rect 1310 354 1506 1132
rect 1672 442 1746 460
rect 210 -248 390 150
rect 782 -248 932 170
rect 210 -310 932 -248
rect 208 -372 932 -310
rect 1312 -208 1518 148
rect 1672 74 1686 442
rect 1730 356 1746 442
rect 1998 356 2244 424
rect 1730 344 2244 356
rect 1730 160 2060 344
rect 1730 74 1746 160
rect 1874 158 2060 160
rect 1998 134 2060 158
rect 2192 134 2244 344
rect 1998 74 2244 134
rect 1672 48 1746 74
rect 208 -794 394 -372
rect 1312 -376 2580 -208
rect 1312 -646 1518 -376
rect 1692 -566 2202 -548
rect 772 -848 1276 -652
rect 772 -1136 982 -848
rect 1324 -1536 1522 -856
rect 1692 -938 1708 -566
rect 1744 -586 2202 -566
rect 1744 -656 2152 -586
rect 1744 -866 1870 -656
rect 1998 -866 2152 -656
rect 1744 -938 2152 -866
rect 1692 -958 2152 -938
rect 2188 -958 2202 -586
rect 2376 -668 2578 -376
rect 2620 -876 3264 -676
rect 1692 -972 2202 -958
rect 2374 -1526 2566 -884
<< via1 >>
rect 214 688 380 932
rect 2060 134 2192 344
rect 1870 -866 1998 -656
<< metal2 >>
rect 202 932 2204 966
rect 202 836 214 932
rect 200 688 214 836
rect 380 842 2204 932
rect 380 688 388 842
rect 200 682 388 688
rect 2018 426 2204 842
rect 1994 344 2242 426
rect 1994 134 2060 344
rect 2192 134 2242 344
rect 1994 86 2242 134
rect 1816 -98 2242 86
rect 1818 -574 2048 -98
rect 1782 -656 2082 -574
rect 1782 -866 1870 -656
rect 1998 -866 2082 -656
rect 1782 -964 2082 -866
use sky130_fd_pr__pfet_g5v0d10v5_6H9SE5  sky130_fd_pr__pfet_g5v0d10v5_6H9SE5_0
timestamp 1695142129
transform 0 1 302 -1 0 263
box -358 -397 358 397
use sky130_fd_pr__pfet_g5v0d10v5_6H9SE5  sky130_fd_pr__pfet_g5v0d10v5_6H9SE5_1
timestamp 1695142129
transform 0 1 1408 -1 0 255
box -358 -397 358 397
use sky130_fd_pr__pfet_g5v0d10v5_6H9SE5  sky130_fd_pr__pfet_g5v0d10v5_6H9SE5_2
timestamp 1695142129
transform 0 1 2472 -1 0 -773
box -358 -397 358 397
use sky130_fd_pr__pfet_g5v0d10v5_6H9SE5  sky130_fd_pr__pfet_g5v0d10v5_6H9SE5_3
timestamp 1695142129
transform 0 1 1424 -1 0 -753
box -358 -397 358 397
use sky130_fd_pr__res_iso_pw_25QSVZ  sky130_fd_pr__res_iso_pw_25QSVZ_0
timestamp 1695142129
transform 1 0 2264 0 1 7507
box -1248 -6017 1248 6017
<< labels >>
rlabel metal1 226 -772 364 -598 1 iin
port 6 n
rlabel metal1 1214 13938 1570 14364 1 vdd
port 1 n
rlabel metal1 1352 -1514 1482 -1302 1 iout
port 4 n
rlabel metal1 2404 -1506 2534 -1294 1 iout_neg
port 3 n
rlabel metal1 3084 -862 3244 -698 1 vbias
port 2 n
rlabel metal1 792 -1108 952 -944 1 vsw
port 5 n
<< end >>
