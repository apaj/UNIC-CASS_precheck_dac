magic
tech sky130A
timestamp 1628284015
<< end >>
