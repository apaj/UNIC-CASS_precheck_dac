magic
tech sky130A
magscale 1 2
timestamp 1697620687
<< viali >>
rect 10842 2674 10884 2884
rect 10860 2166 10898 2378
rect 10858 1688 10896 1894
rect -2522 1442 -2338 1644
rect 10862 1176 10896 1384
rect -1014 220 -916 326
rect 268 192 412 338
rect -1538 -36 -1164 0
rect -512 -54 -138 -18
rect -1494 -382 -1326 -248
rect -520 -568 -152 -534
rect 588 -578 956 -544
rect -800 -926 -680 -782
rect 314 -942 438 -794
<< metal1 >>
rect 10838 2900 10924 2902
rect 10826 2884 10924 2900
rect -1728 2676 -1276 2856
rect -3902 2442 -1276 2676
rect -3902 2436 -3702 2442
rect -3130 2378 -1276 2442
rect -3130 376 -2782 2378
rect -1728 2192 -1276 2378
rect -1708 1694 -1272 1868
rect -2590 1644 -1272 1694
rect -2590 1442 -2522 1644
rect -2338 1442 -1272 1644
rect -2590 1396 -1272 1442
rect -1708 1220 -1272 1396
rect 10330 1196 10744 2848
rect 10826 2674 10842 2884
rect 10884 2674 10924 2884
rect 10826 2656 10924 2674
rect 10838 2378 10924 2656
rect 10838 2166 10860 2378
rect 10898 2166 10924 2378
rect 10838 1894 10924 2166
rect 10838 1688 10858 1894
rect 10896 1688 10924 1894
rect 10838 1384 10924 1688
rect 10838 1176 10862 1384
rect 10896 1222 10924 1384
rect 10896 1176 10926 1222
rect 10838 918 10926 1176
rect 10834 780 10928 918
rect -1458 680 -218 770
rect -1458 424 -1248 680
rect -1006 376 -890 680
rect -430 406 -220 680
rect 10792 580 10992 780
rect -3130 198 -1464 376
rect -3118 184 -1464 198
rect -1242 326 -890 376
rect -1242 220 -1014 326
rect -916 220 -890 326
rect -1242 192 -890 220
rect -814 328 -430 364
rect -814 222 -774 328
rect -676 222 -430 328
rect -814 196 -430 222
rect -216 338 424 352
rect -216 192 268 338
rect 412 192 424 338
rect -2132 36 -1886 184
rect -216 176 424 192
rect -2132 0 -132 36
rect -2132 -36 -1538 0
rect -1164 -10 -132 0
rect -1164 -18 -124 -10
rect -1164 -36 -512 -18
rect -2132 -54 -512 -36
rect -138 -54 -124 -18
rect -2132 -68 -124 -54
rect -2132 -70 -128 -68
rect -1548 -76 -128 -70
rect -1518 -248 -1308 -232
rect -1518 -382 -1494 -248
rect -1326 -382 -1308 -248
rect -1518 -696 -1308 -382
rect -470 -516 -242 -76
rect -544 -518 -138 -516
rect -544 -524 964 -518
rect -544 -534 968 -524
rect -544 -568 -520 -534
rect -152 -544 968 -534
rect -152 -568 588 -544
rect -544 -578 588 -568
rect 956 -578 968 -544
rect -544 -584 968 -578
rect -544 -590 -138 -584
rect 574 -596 968 -584
rect -1512 -700 -1312 -696
rect -94 -764 110 -758
rect -812 -782 -448 -764
rect -812 -926 -800 -782
rect -680 -926 -448 -782
rect -812 -942 -448 -926
rect -224 -936 114 -764
rect 300 -794 664 -774
rect -438 -1426 -254 -996
rect -446 -1634 -254 -1426
rect -94 -1492 110 -936
rect 300 -942 314 -794
rect 438 -942 664 -794
rect 300 -952 664 -942
rect 882 -946 1312 -776
rect 686 -1388 854 -1006
rect -86 -1634 106 -1492
rect 662 -1592 854 -1388
rect 1128 -1324 1312 -946
rect 1128 -1478 1324 -1324
rect 1132 -1528 1324 -1478
rect -448 -1834 -248 -1634
rect -86 -1834 118 -1634
rect 660 -1792 860 -1592
rect 1132 -1728 1332 -1528
<< via1 >>
rect -2522 1442 -2338 1644
rect -1014 220 -916 326
rect -774 222 -676 328
rect 268 192 412 338
rect -1494 -382 -1326 -248
rect -800 -926 -680 -782
rect 314 -942 438 -794
<< metal2 >>
rect -2586 1644 -2232 1706
rect -2586 1442 -2522 1644
rect -2338 1442 -2232 1644
rect -2586 952 -2232 1442
rect -2586 946 -1462 952
rect -2586 836 -636 946
rect -2586 834 -1462 836
rect -2586 830 -2232 834
rect -820 392 -636 836
rect -1050 326 -888 358
rect -1050 220 -1014 326
rect -916 220 -888 326
rect -820 328 -638 392
rect -820 306 -774 328
rect -1050 -154 -888 220
rect -814 222 -774 306
rect -676 222 -638 328
rect -814 196 -638 222
rect 234 338 442 352
rect -1518 -248 -888 -154
rect -1518 -382 -1494 -248
rect -1326 -320 -888 -248
rect 234 192 268 338
rect 412 192 442 338
rect -1326 -382 -892 -320
rect 234 -328 442 192
rect -1518 -412 -892 -382
rect -822 -452 444 -328
rect -822 -782 -666 -452
rect -822 -926 -800 -782
rect -680 -926 -666 -782
rect -822 -946 -666 -926
rect 286 -774 442 -452
rect 286 -794 456 -774
rect 286 -942 314 -794
rect 438 -942 456 -794
rect 286 -960 456 -942
use sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0  XM1
timestamp 1697388883
transform 1 0 -1354 0 1 281
box -358 -397 358 397
use sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0  XM2
timestamp 1697388883
transform 1 0 -326 0 1 263
box -358 -397 358 397
use sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0  XM3
timestamp 1697388883
transform 1 0 -336 0 1 -853
box -358 -397 358 397
use sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0  XM4
timestamp 1697388883
transform 1 0 772 0 1 -863
box -358 -397 358 397
use sky130_fd_pr__res_xhigh_po_0p69_MS44J6  XR1
timestamp 1697384985
transform 0 -1 4534 1 0 1279
box -235 -6398 235 6398
use sky130_fd_pr__res_xhigh_po_0p69_MS44J6  XR2
timestamp 1697384985
transform 0 -1 4532 1 0 1791
box -235 -6398 235 6398
use sky130_fd_pr__res_xhigh_po_0p69_MS44J6  XR3
timestamp 1697384985
transform 0 -1 4534 1 0 2271
box -235 -6398 235 6398
use sky130_fd_pr__res_xhigh_po_0p69_MS44J6  XR4
timestamp 1697384985
transform 0 -1 4518 1 0 2777
box -235 -6398 235 6398
<< labels >>
flabel metal1 10792 580 10992 780 0 FreeSans 1280 0 0 0 vgnd
port 1 nsew
flabel metal1 -3902 2436 -3702 2636 0 FreeSans 1280 0 0 0 vsup
port 0 nsew
flabel metal1 -1512 -700 -1312 -500 0 FreeSans 1280 0 0 0 iref
port 2 nsew
flabel metal1 -448 -1834 -248 -1634 0 FreeSans 1280 0 0 0 vsw
port 3 nsew
flabel metal1 -82 -1834 118 -1634 0 FreeSans 1280 0 0 0 iout
port 4 nsew
flabel metal1 1132 -1728 1332 -1528 0 FreeSans 1280 0 0 0 iout_n
port 5 nsew
flabel metal1 660 -1792 860 -1592 0 FreeSans 1280 0 0 0 vbias
port 6 nsew
rlabel metal1 10330 1196 10744 2848 1 parR
rlabel metal2 234 -452 442 192 1 sourceM3M4
rlabel metal2 -2586 834 -1462 952 1 sourceM2
<< end >>
