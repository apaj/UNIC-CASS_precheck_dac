magic
tech sky130A
magscale 1 2
timestamp 1697534501
<< nwell >>
rect -2949 -26297 2949 26297
<< mvpmos >>
rect -2691 -26000 -2591 26000
rect -2413 -26000 -2313 26000
rect -2135 -26000 -2035 26000
rect -1857 -26000 -1757 26000
rect -1579 -26000 -1479 26000
rect -1301 -26000 -1201 26000
rect -1023 -26000 -923 26000
rect -745 -26000 -645 26000
rect -467 -26000 -367 26000
rect -189 -26000 -89 26000
rect 89 -26000 189 26000
rect 367 -26000 467 26000
rect 645 -26000 745 26000
rect 923 -26000 1023 26000
rect 1201 -26000 1301 26000
rect 1479 -26000 1579 26000
rect 1757 -26000 1857 26000
rect 2035 -26000 2135 26000
rect 2313 -26000 2413 26000
rect 2591 -26000 2691 26000
<< mvpdiff >>
rect -2749 25988 -2691 26000
rect -2749 -25988 -2737 25988
rect -2703 -25988 -2691 25988
rect -2749 -26000 -2691 -25988
rect -2591 25988 -2533 26000
rect -2591 -25988 -2579 25988
rect -2545 -25988 -2533 25988
rect -2591 -26000 -2533 -25988
rect -2471 25988 -2413 26000
rect -2471 -25988 -2459 25988
rect -2425 -25988 -2413 25988
rect -2471 -26000 -2413 -25988
rect -2313 25988 -2255 26000
rect -2313 -25988 -2301 25988
rect -2267 -25988 -2255 25988
rect -2313 -26000 -2255 -25988
rect -2193 25988 -2135 26000
rect -2193 -25988 -2181 25988
rect -2147 -25988 -2135 25988
rect -2193 -26000 -2135 -25988
rect -2035 25988 -1977 26000
rect -2035 -25988 -2023 25988
rect -1989 -25988 -1977 25988
rect -2035 -26000 -1977 -25988
rect -1915 25988 -1857 26000
rect -1915 -25988 -1903 25988
rect -1869 -25988 -1857 25988
rect -1915 -26000 -1857 -25988
rect -1757 25988 -1699 26000
rect -1757 -25988 -1745 25988
rect -1711 -25988 -1699 25988
rect -1757 -26000 -1699 -25988
rect -1637 25988 -1579 26000
rect -1637 -25988 -1625 25988
rect -1591 -25988 -1579 25988
rect -1637 -26000 -1579 -25988
rect -1479 25988 -1421 26000
rect -1479 -25988 -1467 25988
rect -1433 -25988 -1421 25988
rect -1479 -26000 -1421 -25988
rect -1359 25988 -1301 26000
rect -1359 -25988 -1347 25988
rect -1313 -25988 -1301 25988
rect -1359 -26000 -1301 -25988
rect -1201 25988 -1143 26000
rect -1201 -25988 -1189 25988
rect -1155 -25988 -1143 25988
rect -1201 -26000 -1143 -25988
rect -1081 25988 -1023 26000
rect -1081 -25988 -1069 25988
rect -1035 -25988 -1023 25988
rect -1081 -26000 -1023 -25988
rect -923 25988 -865 26000
rect -923 -25988 -911 25988
rect -877 -25988 -865 25988
rect -923 -26000 -865 -25988
rect -803 25988 -745 26000
rect -803 -25988 -791 25988
rect -757 -25988 -745 25988
rect -803 -26000 -745 -25988
rect -645 25988 -587 26000
rect -645 -25988 -633 25988
rect -599 -25988 -587 25988
rect -645 -26000 -587 -25988
rect -525 25988 -467 26000
rect -525 -25988 -513 25988
rect -479 -25988 -467 25988
rect -525 -26000 -467 -25988
rect -367 25988 -309 26000
rect -367 -25988 -355 25988
rect -321 -25988 -309 25988
rect -367 -26000 -309 -25988
rect -247 25988 -189 26000
rect -247 -25988 -235 25988
rect -201 -25988 -189 25988
rect -247 -26000 -189 -25988
rect -89 25988 -31 26000
rect -89 -25988 -77 25988
rect -43 -25988 -31 25988
rect -89 -26000 -31 -25988
rect 31 25988 89 26000
rect 31 -25988 43 25988
rect 77 -25988 89 25988
rect 31 -26000 89 -25988
rect 189 25988 247 26000
rect 189 -25988 201 25988
rect 235 -25988 247 25988
rect 189 -26000 247 -25988
rect 309 25988 367 26000
rect 309 -25988 321 25988
rect 355 -25988 367 25988
rect 309 -26000 367 -25988
rect 467 25988 525 26000
rect 467 -25988 479 25988
rect 513 -25988 525 25988
rect 467 -26000 525 -25988
rect 587 25988 645 26000
rect 587 -25988 599 25988
rect 633 -25988 645 25988
rect 587 -26000 645 -25988
rect 745 25988 803 26000
rect 745 -25988 757 25988
rect 791 -25988 803 25988
rect 745 -26000 803 -25988
rect 865 25988 923 26000
rect 865 -25988 877 25988
rect 911 -25988 923 25988
rect 865 -26000 923 -25988
rect 1023 25988 1081 26000
rect 1023 -25988 1035 25988
rect 1069 -25988 1081 25988
rect 1023 -26000 1081 -25988
rect 1143 25988 1201 26000
rect 1143 -25988 1155 25988
rect 1189 -25988 1201 25988
rect 1143 -26000 1201 -25988
rect 1301 25988 1359 26000
rect 1301 -25988 1313 25988
rect 1347 -25988 1359 25988
rect 1301 -26000 1359 -25988
rect 1421 25988 1479 26000
rect 1421 -25988 1433 25988
rect 1467 -25988 1479 25988
rect 1421 -26000 1479 -25988
rect 1579 25988 1637 26000
rect 1579 -25988 1591 25988
rect 1625 -25988 1637 25988
rect 1579 -26000 1637 -25988
rect 1699 25988 1757 26000
rect 1699 -25988 1711 25988
rect 1745 -25988 1757 25988
rect 1699 -26000 1757 -25988
rect 1857 25988 1915 26000
rect 1857 -25988 1869 25988
rect 1903 -25988 1915 25988
rect 1857 -26000 1915 -25988
rect 1977 25988 2035 26000
rect 1977 -25988 1989 25988
rect 2023 -25988 2035 25988
rect 1977 -26000 2035 -25988
rect 2135 25988 2193 26000
rect 2135 -25988 2147 25988
rect 2181 -25988 2193 25988
rect 2135 -26000 2193 -25988
rect 2255 25988 2313 26000
rect 2255 -25988 2267 25988
rect 2301 -25988 2313 25988
rect 2255 -26000 2313 -25988
rect 2413 25988 2471 26000
rect 2413 -25988 2425 25988
rect 2459 -25988 2471 25988
rect 2413 -26000 2471 -25988
rect 2533 25988 2591 26000
rect 2533 -25988 2545 25988
rect 2579 -25988 2591 25988
rect 2533 -26000 2591 -25988
rect 2691 25988 2749 26000
rect 2691 -25988 2703 25988
rect 2737 -25988 2749 25988
rect 2691 -26000 2749 -25988
<< mvpdiffc >>
rect -2737 -25988 -2703 25988
rect -2579 -25988 -2545 25988
rect -2459 -25988 -2425 25988
rect -2301 -25988 -2267 25988
rect -2181 -25988 -2147 25988
rect -2023 -25988 -1989 25988
rect -1903 -25988 -1869 25988
rect -1745 -25988 -1711 25988
rect -1625 -25988 -1591 25988
rect -1467 -25988 -1433 25988
rect -1347 -25988 -1313 25988
rect -1189 -25988 -1155 25988
rect -1069 -25988 -1035 25988
rect -911 -25988 -877 25988
rect -791 -25988 -757 25988
rect -633 -25988 -599 25988
rect -513 -25988 -479 25988
rect -355 -25988 -321 25988
rect -235 -25988 -201 25988
rect -77 -25988 -43 25988
rect 43 -25988 77 25988
rect 201 -25988 235 25988
rect 321 -25988 355 25988
rect 479 -25988 513 25988
rect 599 -25988 633 25988
rect 757 -25988 791 25988
rect 877 -25988 911 25988
rect 1035 -25988 1069 25988
rect 1155 -25988 1189 25988
rect 1313 -25988 1347 25988
rect 1433 -25988 1467 25988
rect 1591 -25988 1625 25988
rect 1711 -25988 1745 25988
rect 1869 -25988 1903 25988
rect 1989 -25988 2023 25988
rect 2147 -25988 2181 25988
rect 2267 -25988 2301 25988
rect 2425 -25988 2459 25988
rect 2545 -25988 2579 25988
rect 2703 -25988 2737 25988
<< mvnsubdiff >>
rect -2883 26219 2883 26231
rect -2883 26185 -2775 26219
rect 2775 26185 2883 26219
rect -2883 26173 2883 26185
rect -2883 26123 -2825 26173
rect -2883 -26123 -2871 26123
rect -2837 -26123 -2825 26123
rect 2825 26123 2883 26173
rect -2883 -26173 -2825 -26123
rect 2825 -26123 2837 26123
rect 2871 -26123 2883 26123
rect 2825 -26173 2883 -26123
rect -2883 -26185 2883 -26173
rect -2883 -26219 -2775 -26185
rect 2775 -26219 2883 -26185
rect -2883 -26231 2883 -26219
<< mvnsubdiffcont >>
rect -2775 26185 2775 26219
rect -2871 -26123 -2837 26123
rect 2837 -26123 2871 26123
rect -2775 -26219 2775 -26185
<< poly >>
rect -2691 26081 -2591 26097
rect -2691 26047 -2675 26081
rect -2607 26047 -2591 26081
rect -2691 26000 -2591 26047
rect -2413 26081 -2313 26097
rect -2413 26047 -2397 26081
rect -2329 26047 -2313 26081
rect -2413 26000 -2313 26047
rect -2135 26081 -2035 26097
rect -2135 26047 -2119 26081
rect -2051 26047 -2035 26081
rect -2135 26000 -2035 26047
rect -1857 26081 -1757 26097
rect -1857 26047 -1841 26081
rect -1773 26047 -1757 26081
rect -1857 26000 -1757 26047
rect -1579 26081 -1479 26097
rect -1579 26047 -1563 26081
rect -1495 26047 -1479 26081
rect -1579 26000 -1479 26047
rect -1301 26081 -1201 26097
rect -1301 26047 -1285 26081
rect -1217 26047 -1201 26081
rect -1301 26000 -1201 26047
rect -1023 26081 -923 26097
rect -1023 26047 -1007 26081
rect -939 26047 -923 26081
rect -1023 26000 -923 26047
rect -745 26081 -645 26097
rect -745 26047 -729 26081
rect -661 26047 -645 26081
rect -745 26000 -645 26047
rect -467 26081 -367 26097
rect -467 26047 -451 26081
rect -383 26047 -367 26081
rect -467 26000 -367 26047
rect -189 26081 -89 26097
rect -189 26047 -173 26081
rect -105 26047 -89 26081
rect -189 26000 -89 26047
rect 89 26081 189 26097
rect 89 26047 105 26081
rect 173 26047 189 26081
rect 89 26000 189 26047
rect 367 26081 467 26097
rect 367 26047 383 26081
rect 451 26047 467 26081
rect 367 26000 467 26047
rect 645 26081 745 26097
rect 645 26047 661 26081
rect 729 26047 745 26081
rect 645 26000 745 26047
rect 923 26081 1023 26097
rect 923 26047 939 26081
rect 1007 26047 1023 26081
rect 923 26000 1023 26047
rect 1201 26081 1301 26097
rect 1201 26047 1217 26081
rect 1285 26047 1301 26081
rect 1201 26000 1301 26047
rect 1479 26081 1579 26097
rect 1479 26047 1495 26081
rect 1563 26047 1579 26081
rect 1479 26000 1579 26047
rect 1757 26081 1857 26097
rect 1757 26047 1773 26081
rect 1841 26047 1857 26081
rect 1757 26000 1857 26047
rect 2035 26081 2135 26097
rect 2035 26047 2051 26081
rect 2119 26047 2135 26081
rect 2035 26000 2135 26047
rect 2313 26081 2413 26097
rect 2313 26047 2329 26081
rect 2397 26047 2413 26081
rect 2313 26000 2413 26047
rect 2591 26081 2691 26097
rect 2591 26047 2607 26081
rect 2675 26047 2691 26081
rect 2591 26000 2691 26047
rect -2691 -26047 -2591 -26000
rect -2691 -26081 -2675 -26047
rect -2607 -26081 -2591 -26047
rect -2691 -26097 -2591 -26081
rect -2413 -26047 -2313 -26000
rect -2413 -26081 -2397 -26047
rect -2329 -26081 -2313 -26047
rect -2413 -26097 -2313 -26081
rect -2135 -26047 -2035 -26000
rect -2135 -26081 -2119 -26047
rect -2051 -26081 -2035 -26047
rect -2135 -26097 -2035 -26081
rect -1857 -26047 -1757 -26000
rect -1857 -26081 -1841 -26047
rect -1773 -26081 -1757 -26047
rect -1857 -26097 -1757 -26081
rect -1579 -26047 -1479 -26000
rect -1579 -26081 -1563 -26047
rect -1495 -26081 -1479 -26047
rect -1579 -26097 -1479 -26081
rect -1301 -26047 -1201 -26000
rect -1301 -26081 -1285 -26047
rect -1217 -26081 -1201 -26047
rect -1301 -26097 -1201 -26081
rect -1023 -26047 -923 -26000
rect -1023 -26081 -1007 -26047
rect -939 -26081 -923 -26047
rect -1023 -26097 -923 -26081
rect -745 -26047 -645 -26000
rect -745 -26081 -729 -26047
rect -661 -26081 -645 -26047
rect -745 -26097 -645 -26081
rect -467 -26047 -367 -26000
rect -467 -26081 -451 -26047
rect -383 -26081 -367 -26047
rect -467 -26097 -367 -26081
rect -189 -26047 -89 -26000
rect -189 -26081 -173 -26047
rect -105 -26081 -89 -26047
rect -189 -26097 -89 -26081
rect 89 -26047 189 -26000
rect 89 -26081 105 -26047
rect 173 -26081 189 -26047
rect 89 -26097 189 -26081
rect 367 -26047 467 -26000
rect 367 -26081 383 -26047
rect 451 -26081 467 -26047
rect 367 -26097 467 -26081
rect 645 -26047 745 -26000
rect 645 -26081 661 -26047
rect 729 -26081 745 -26047
rect 645 -26097 745 -26081
rect 923 -26047 1023 -26000
rect 923 -26081 939 -26047
rect 1007 -26081 1023 -26047
rect 923 -26097 1023 -26081
rect 1201 -26047 1301 -26000
rect 1201 -26081 1217 -26047
rect 1285 -26081 1301 -26047
rect 1201 -26097 1301 -26081
rect 1479 -26047 1579 -26000
rect 1479 -26081 1495 -26047
rect 1563 -26081 1579 -26047
rect 1479 -26097 1579 -26081
rect 1757 -26047 1857 -26000
rect 1757 -26081 1773 -26047
rect 1841 -26081 1857 -26047
rect 1757 -26097 1857 -26081
rect 2035 -26047 2135 -26000
rect 2035 -26081 2051 -26047
rect 2119 -26081 2135 -26047
rect 2035 -26097 2135 -26081
rect 2313 -26047 2413 -26000
rect 2313 -26081 2329 -26047
rect 2397 -26081 2413 -26047
rect 2313 -26097 2413 -26081
rect 2591 -26047 2691 -26000
rect 2591 -26081 2607 -26047
rect 2675 -26081 2691 -26047
rect 2591 -26097 2691 -26081
<< polycont >>
rect -2675 26047 -2607 26081
rect -2397 26047 -2329 26081
rect -2119 26047 -2051 26081
rect -1841 26047 -1773 26081
rect -1563 26047 -1495 26081
rect -1285 26047 -1217 26081
rect -1007 26047 -939 26081
rect -729 26047 -661 26081
rect -451 26047 -383 26081
rect -173 26047 -105 26081
rect 105 26047 173 26081
rect 383 26047 451 26081
rect 661 26047 729 26081
rect 939 26047 1007 26081
rect 1217 26047 1285 26081
rect 1495 26047 1563 26081
rect 1773 26047 1841 26081
rect 2051 26047 2119 26081
rect 2329 26047 2397 26081
rect 2607 26047 2675 26081
rect -2675 -26081 -2607 -26047
rect -2397 -26081 -2329 -26047
rect -2119 -26081 -2051 -26047
rect -1841 -26081 -1773 -26047
rect -1563 -26081 -1495 -26047
rect -1285 -26081 -1217 -26047
rect -1007 -26081 -939 -26047
rect -729 -26081 -661 -26047
rect -451 -26081 -383 -26047
rect -173 -26081 -105 -26047
rect 105 -26081 173 -26047
rect 383 -26081 451 -26047
rect 661 -26081 729 -26047
rect 939 -26081 1007 -26047
rect 1217 -26081 1285 -26047
rect 1495 -26081 1563 -26047
rect 1773 -26081 1841 -26047
rect 2051 -26081 2119 -26047
rect 2329 -26081 2397 -26047
rect 2607 -26081 2675 -26047
<< locali >>
rect -2871 26185 -2775 26219
rect 2775 26185 2871 26219
rect -2871 26123 -2837 26185
rect 2837 26123 2871 26185
rect -2691 26047 -2675 26081
rect -2607 26047 -2591 26081
rect -2413 26047 -2397 26081
rect -2329 26047 -2313 26081
rect -2135 26047 -2119 26081
rect -2051 26047 -2035 26081
rect -1857 26047 -1841 26081
rect -1773 26047 -1757 26081
rect -1579 26047 -1563 26081
rect -1495 26047 -1479 26081
rect -1301 26047 -1285 26081
rect -1217 26047 -1201 26081
rect -1023 26047 -1007 26081
rect -939 26047 -923 26081
rect -745 26047 -729 26081
rect -661 26047 -645 26081
rect -467 26047 -451 26081
rect -383 26047 -367 26081
rect -189 26047 -173 26081
rect -105 26047 -89 26081
rect 89 26047 105 26081
rect 173 26047 189 26081
rect 367 26047 383 26081
rect 451 26047 467 26081
rect 645 26047 661 26081
rect 729 26047 745 26081
rect 923 26047 939 26081
rect 1007 26047 1023 26081
rect 1201 26047 1217 26081
rect 1285 26047 1301 26081
rect 1479 26047 1495 26081
rect 1563 26047 1579 26081
rect 1757 26047 1773 26081
rect 1841 26047 1857 26081
rect 2035 26047 2051 26081
rect 2119 26047 2135 26081
rect 2313 26047 2329 26081
rect 2397 26047 2413 26081
rect 2591 26047 2607 26081
rect 2675 26047 2691 26081
rect -2737 25988 -2703 26004
rect -2737 -26004 -2703 -25988
rect -2579 25988 -2545 26004
rect -2579 -26004 -2545 -25988
rect -2459 25988 -2425 26004
rect -2459 -26004 -2425 -25988
rect -2301 25988 -2267 26004
rect -2301 -26004 -2267 -25988
rect -2181 25988 -2147 26004
rect -2181 -26004 -2147 -25988
rect -2023 25988 -1989 26004
rect -2023 -26004 -1989 -25988
rect -1903 25988 -1869 26004
rect -1903 -26004 -1869 -25988
rect -1745 25988 -1711 26004
rect -1745 -26004 -1711 -25988
rect -1625 25988 -1591 26004
rect -1625 -26004 -1591 -25988
rect -1467 25988 -1433 26004
rect -1467 -26004 -1433 -25988
rect -1347 25988 -1313 26004
rect -1347 -26004 -1313 -25988
rect -1189 25988 -1155 26004
rect -1189 -26004 -1155 -25988
rect -1069 25988 -1035 26004
rect -1069 -26004 -1035 -25988
rect -911 25988 -877 26004
rect -911 -26004 -877 -25988
rect -791 25988 -757 26004
rect -791 -26004 -757 -25988
rect -633 25988 -599 26004
rect -633 -26004 -599 -25988
rect -513 25988 -479 26004
rect -513 -26004 -479 -25988
rect -355 25988 -321 26004
rect -355 -26004 -321 -25988
rect -235 25988 -201 26004
rect -235 -26004 -201 -25988
rect -77 25988 -43 26004
rect -77 -26004 -43 -25988
rect 43 25988 77 26004
rect 43 -26004 77 -25988
rect 201 25988 235 26004
rect 201 -26004 235 -25988
rect 321 25988 355 26004
rect 321 -26004 355 -25988
rect 479 25988 513 26004
rect 479 -26004 513 -25988
rect 599 25988 633 26004
rect 599 -26004 633 -25988
rect 757 25988 791 26004
rect 757 -26004 791 -25988
rect 877 25988 911 26004
rect 877 -26004 911 -25988
rect 1035 25988 1069 26004
rect 1035 -26004 1069 -25988
rect 1155 25988 1189 26004
rect 1155 -26004 1189 -25988
rect 1313 25988 1347 26004
rect 1313 -26004 1347 -25988
rect 1433 25988 1467 26004
rect 1433 -26004 1467 -25988
rect 1591 25988 1625 26004
rect 1591 -26004 1625 -25988
rect 1711 25988 1745 26004
rect 1711 -26004 1745 -25988
rect 1869 25988 1903 26004
rect 1869 -26004 1903 -25988
rect 1989 25988 2023 26004
rect 1989 -26004 2023 -25988
rect 2147 25988 2181 26004
rect 2147 -26004 2181 -25988
rect 2267 25988 2301 26004
rect 2267 -26004 2301 -25988
rect 2425 25988 2459 26004
rect 2425 -26004 2459 -25988
rect 2545 25988 2579 26004
rect 2545 -26004 2579 -25988
rect 2703 25988 2737 26004
rect 2703 -26004 2737 -25988
rect -2691 -26081 -2675 -26047
rect -2607 -26081 -2591 -26047
rect -2413 -26081 -2397 -26047
rect -2329 -26081 -2313 -26047
rect -2135 -26081 -2119 -26047
rect -2051 -26081 -2035 -26047
rect -1857 -26081 -1841 -26047
rect -1773 -26081 -1757 -26047
rect -1579 -26081 -1563 -26047
rect -1495 -26081 -1479 -26047
rect -1301 -26081 -1285 -26047
rect -1217 -26081 -1201 -26047
rect -1023 -26081 -1007 -26047
rect -939 -26081 -923 -26047
rect -745 -26081 -729 -26047
rect -661 -26081 -645 -26047
rect -467 -26081 -451 -26047
rect -383 -26081 -367 -26047
rect -189 -26081 -173 -26047
rect -105 -26081 -89 -26047
rect 89 -26081 105 -26047
rect 173 -26081 189 -26047
rect 367 -26081 383 -26047
rect 451 -26081 467 -26047
rect 645 -26081 661 -26047
rect 729 -26081 745 -26047
rect 923 -26081 939 -26047
rect 1007 -26081 1023 -26047
rect 1201 -26081 1217 -26047
rect 1285 -26081 1301 -26047
rect 1479 -26081 1495 -26047
rect 1563 -26081 1579 -26047
rect 1757 -26081 1773 -26047
rect 1841 -26081 1857 -26047
rect 2035 -26081 2051 -26047
rect 2119 -26081 2135 -26047
rect 2313 -26081 2329 -26047
rect 2397 -26081 2413 -26047
rect 2591 -26081 2607 -26047
rect 2675 -26081 2691 -26047
rect -2871 -26185 -2837 -26123
rect 2837 -26185 2871 -26123
rect -2871 -26219 -2775 -26185
rect 2775 -26219 2871 -26185
<< viali >>
rect -2675 26047 -2607 26081
rect -2397 26047 -2329 26081
rect -2119 26047 -2051 26081
rect -1841 26047 -1773 26081
rect -1563 26047 -1495 26081
rect -1285 26047 -1217 26081
rect -1007 26047 -939 26081
rect -729 26047 -661 26081
rect -451 26047 -383 26081
rect -173 26047 -105 26081
rect 105 26047 173 26081
rect 383 26047 451 26081
rect 661 26047 729 26081
rect 939 26047 1007 26081
rect 1217 26047 1285 26081
rect 1495 26047 1563 26081
rect 1773 26047 1841 26081
rect 2051 26047 2119 26081
rect 2329 26047 2397 26081
rect 2607 26047 2675 26081
rect -2737 -25988 -2703 25988
rect -2579 -25988 -2545 25988
rect -2459 -25988 -2425 25988
rect -2301 -25988 -2267 25988
rect -2181 -25988 -2147 25988
rect -2023 -25988 -1989 25988
rect -1903 -25988 -1869 25988
rect -1745 -25988 -1711 25988
rect -1625 -25988 -1591 25988
rect -1467 -25988 -1433 25988
rect -1347 -25988 -1313 25988
rect -1189 -25988 -1155 25988
rect -1069 -25988 -1035 25988
rect -911 -25988 -877 25988
rect -791 -25988 -757 25988
rect -633 -25988 -599 25988
rect -513 -25988 -479 25988
rect -355 -25988 -321 25988
rect -235 -25988 -201 25988
rect -77 -25988 -43 25988
rect 43 -25988 77 25988
rect 201 -25988 235 25988
rect 321 -25988 355 25988
rect 479 -25988 513 25988
rect 599 -25988 633 25988
rect 757 -25988 791 25988
rect 877 -25988 911 25988
rect 1035 -25988 1069 25988
rect 1155 -25988 1189 25988
rect 1313 -25988 1347 25988
rect 1433 -25988 1467 25988
rect 1591 -25988 1625 25988
rect 1711 -25988 1745 25988
rect 1869 -25988 1903 25988
rect 1989 -25988 2023 25988
rect 2147 -25988 2181 25988
rect 2267 -25988 2301 25988
rect 2425 -25988 2459 25988
rect 2545 -25988 2579 25988
rect 2703 -25988 2737 25988
rect -2675 -26081 -2607 -26047
rect -2397 -26081 -2329 -26047
rect -2119 -26081 -2051 -26047
rect -1841 -26081 -1773 -26047
rect -1563 -26081 -1495 -26047
rect -1285 -26081 -1217 -26047
rect -1007 -26081 -939 -26047
rect -729 -26081 -661 -26047
rect -451 -26081 -383 -26047
rect -173 -26081 -105 -26047
rect 105 -26081 173 -26047
rect 383 -26081 451 -26047
rect 661 -26081 729 -26047
rect 939 -26081 1007 -26047
rect 1217 -26081 1285 -26047
rect 1495 -26081 1563 -26047
rect 1773 -26081 1841 -26047
rect 2051 -26081 2119 -26047
rect 2329 -26081 2397 -26047
rect 2607 -26081 2675 -26047
<< metal1 >>
rect -2687 26081 -2595 26087
rect -2687 26047 -2675 26081
rect -2607 26047 -2595 26081
rect -2687 26041 -2595 26047
rect -2409 26081 -2317 26087
rect -2409 26047 -2397 26081
rect -2329 26047 -2317 26081
rect -2409 26041 -2317 26047
rect -2131 26081 -2039 26087
rect -2131 26047 -2119 26081
rect -2051 26047 -2039 26081
rect -2131 26041 -2039 26047
rect -1853 26081 -1761 26087
rect -1853 26047 -1841 26081
rect -1773 26047 -1761 26081
rect -1853 26041 -1761 26047
rect -1575 26081 -1483 26087
rect -1575 26047 -1563 26081
rect -1495 26047 -1483 26081
rect -1575 26041 -1483 26047
rect -1297 26081 -1205 26087
rect -1297 26047 -1285 26081
rect -1217 26047 -1205 26081
rect -1297 26041 -1205 26047
rect -1019 26081 -927 26087
rect -1019 26047 -1007 26081
rect -939 26047 -927 26081
rect -1019 26041 -927 26047
rect -741 26081 -649 26087
rect -741 26047 -729 26081
rect -661 26047 -649 26081
rect -741 26041 -649 26047
rect -463 26081 -371 26087
rect -463 26047 -451 26081
rect -383 26047 -371 26081
rect -463 26041 -371 26047
rect -185 26081 -93 26087
rect -185 26047 -173 26081
rect -105 26047 -93 26081
rect -185 26041 -93 26047
rect 93 26081 185 26087
rect 93 26047 105 26081
rect 173 26047 185 26081
rect 93 26041 185 26047
rect 371 26081 463 26087
rect 371 26047 383 26081
rect 451 26047 463 26081
rect 371 26041 463 26047
rect 649 26081 741 26087
rect 649 26047 661 26081
rect 729 26047 741 26081
rect 649 26041 741 26047
rect 927 26081 1019 26087
rect 927 26047 939 26081
rect 1007 26047 1019 26081
rect 927 26041 1019 26047
rect 1205 26081 1297 26087
rect 1205 26047 1217 26081
rect 1285 26047 1297 26081
rect 1205 26041 1297 26047
rect 1483 26081 1575 26087
rect 1483 26047 1495 26081
rect 1563 26047 1575 26081
rect 1483 26041 1575 26047
rect 1761 26081 1853 26087
rect 1761 26047 1773 26081
rect 1841 26047 1853 26081
rect 1761 26041 1853 26047
rect 2039 26081 2131 26087
rect 2039 26047 2051 26081
rect 2119 26047 2131 26081
rect 2039 26041 2131 26047
rect 2317 26081 2409 26087
rect 2317 26047 2329 26081
rect 2397 26047 2409 26081
rect 2317 26041 2409 26047
rect 2595 26081 2687 26087
rect 2595 26047 2607 26081
rect 2675 26047 2687 26081
rect 2595 26041 2687 26047
rect -2743 25988 -2697 26000
rect -2743 -25988 -2737 25988
rect -2703 -25988 -2697 25988
rect -2743 -26000 -2697 -25988
rect -2585 25988 -2539 26000
rect -2585 -25988 -2579 25988
rect -2545 -25988 -2539 25988
rect -2585 -26000 -2539 -25988
rect -2465 25988 -2419 26000
rect -2465 -25988 -2459 25988
rect -2425 -25988 -2419 25988
rect -2465 -26000 -2419 -25988
rect -2307 25988 -2261 26000
rect -2307 -25988 -2301 25988
rect -2267 -25988 -2261 25988
rect -2307 -26000 -2261 -25988
rect -2187 25988 -2141 26000
rect -2187 -25988 -2181 25988
rect -2147 -25988 -2141 25988
rect -2187 -26000 -2141 -25988
rect -2029 25988 -1983 26000
rect -2029 -25988 -2023 25988
rect -1989 -25988 -1983 25988
rect -2029 -26000 -1983 -25988
rect -1909 25988 -1863 26000
rect -1909 -25988 -1903 25988
rect -1869 -25988 -1863 25988
rect -1909 -26000 -1863 -25988
rect -1751 25988 -1705 26000
rect -1751 -25988 -1745 25988
rect -1711 -25988 -1705 25988
rect -1751 -26000 -1705 -25988
rect -1631 25988 -1585 26000
rect -1631 -25988 -1625 25988
rect -1591 -25988 -1585 25988
rect -1631 -26000 -1585 -25988
rect -1473 25988 -1427 26000
rect -1473 -25988 -1467 25988
rect -1433 -25988 -1427 25988
rect -1473 -26000 -1427 -25988
rect -1353 25988 -1307 26000
rect -1353 -25988 -1347 25988
rect -1313 -25988 -1307 25988
rect -1353 -26000 -1307 -25988
rect -1195 25988 -1149 26000
rect -1195 -25988 -1189 25988
rect -1155 -25988 -1149 25988
rect -1195 -26000 -1149 -25988
rect -1075 25988 -1029 26000
rect -1075 -25988 -1069 25988
rect -1035 -25988 -1029 25988
rect -1075 -26000 -1029 -25988
rect -917 25988 -871 26000
rect -917 -25988 -911 25988
rect -877 -25988 -871 25988
rect -917 -26000 -871 -25988
rect -797 25988 -751 26000
rect -797 -25988 -791 25988
rect -757 -25988 -751 25988
rect -797 -26000 -751 -25988
rect -639 25988 -593 26000
rect -639 -25988 -633 25988
rect -599 -25988 -593 25988
rect -639 -26000 -593 -25988
rect -519 25988 -473 26000
rect -519 -25988 -513 25988
rect -479 -25988 -473 25988
rect -519 -26000 -473 -25988
rect -361 25988 -315 26000
rect -361 -25988 -355 25988
rect -321 -25988 -315 25988
rect -361 -26000 -315 -25988
rect -241 25988 -195 26000
rect -241 -25988 -235 25988
rect -201 -25988 -195 25988
rect -241 -26000 -195 -25988
rect -83 25988 -37 26000
rect -83 -25988 -77 25988
rect -43 -25988 -37 25988
rect -83 -26000 -37 -25988
rect 37 25988 83 26000
rect 37 -25988 43 25988
rect 77 -25988 83 25988
rect 37 -26000 83 -25988
rect 195 25988 241 26000
rect 195 -25988 201 25988
rect 235 -25988 241 25988
rect 195 -26000 241 -25988
rect 315 25988 361 26000
rect 315 -25988 321 25988
rect 355 -25988 361 25988
rect 315 -26000 361 -25988
rect 473 25988 519 26000
rect 473 -25988 479 25988
rect 513 -25988 519 25988
rect 473 -26000 519 -25988
rect 593 25988 639 26000
rect 593 -25988 599 25988
rect 633 -25988 639 25988
rect 593 -26000 639 -25988
rect 751 25988 797 26000
rect 751 -25988 757 25988
rect 791 -25988 797 25988
rect 751 -26000 797 -25988
rect 871 25988 917 26000
rect 871 -25988 877 25988
rect 911 -25988 917 25988
rect 871 -26000 917 -25988
rect 1029 25988 1075 26000
rect 1029 -25988 1035 25988
rect 1069 -25988 1075 25988
rect 1029 -26000 1075 -25988
rect 1149 25988 1195 26000
rect 1149 -25988 1155 25988
rect 1189 -25988 1195 25988
rect 1149 -26000 1195 -25988
rect 1307 25988 1353 26000
rect 1307 -25988 1313 25988
rect 1347 -25988 1353 25988
rect 1307 -26000 1353 -25988
rect 1427 25988 1473 26000
rect 1427 -25988 1433 25988
rect 1467 -25988 1473 25988
rect 1427 -26000 1473 -25988
rect 1585 25988 1631 26000
rect 1585 -25988 1591 25988
rect 1625 -25988 1631 25988
rect 1585 -26000 1631 -25988
rect 1705 25988 1751 26000
rect 1705 -25988 1711 25988
rect 1745 -25988 1751 25988
rect 1705 -26000 1751 -25988
rect 1863 25988 1909 26000
rect 1863 -25988 1869 25988
rect 1903 -25988 1909 25988
rect 1863 -26000 1909 -25988
rect 1983 25988 2029 26000
rect 1983 -25988 1989 25988
rect 2023 -25988 2029 25988
rect 1983 -26000 2029 -25988
rect 2141 25988 2187 26000
rect 2141 -25988 2147 25988
rect 2181 -25988 2187 25988
rect 2141 -26000 2187 -25988
rect 2261 25988 2307 26000
rect 2261 -25988 2267 25988
rect 2301 -25988 2307 25988
rect 2261 -26000 2307 -25988
rect 2419 25988 2465 26000
rect 2419 -25988 2425 25988
rect 2459 -25988 2465 25988
rect 2419 -26000 2465 -25988
rect 2539 25988 2585 26000
rect 2539 -25988 2545 25988
rect 2579 -25988 2585 25988
rect 2539 -26000 2585 -25988
rect 2697 25988 2743 26000
rect 2697 -25988 2703 25988
rect 2737 -25988 2743 25988
rect 2697 -26000 2743 -25988
rect -2687 -26047 -2595 -26041
rect -2687 -26081 -2675 -26047
rect -2607 -26081 -2595 -26047
rect -2687 -26087 -2595 -26081
rect -2409 -26047 -2317 -26041
rect -2409 -26081 -2397 -26047
rect -2329 -26081 -2317 -26047
rect -2409 -26087 -2317 -26081
rect -2131 -26047 -2039 -26041
rect -2131 -26081 -2119 -26047
rect -2051 -26081 -2039 -26047
rect -2131 -26087 -2039 -26081
rect -1853 -26047 -1761 -26041
rect -1853 -26081 -1841 -26047
rect -1773 -26081 -1761 -26047
rect -1853 -26087 -1761 -26081
rect -1575 -26047 -1483 -26041
rect -1575 -26081 -1563 -26047
rect -1495 -26081 -1483 -26047
rect -1575 -26087 -1483 -26081
rect -1297 -26047 -1205 -26041
rect -1297 -26081 -1285 -26047
rect -1217 -26081 -1205 -26047
rect -1297 -26087 -1205 -26081
rect -1019 -26047 -927 -26041
rect -1019 -26081 -1007 -26047
rect -939 -26081 -927 -26047
rect -1019 -26087 -927 -26081
rect -741 -26047 -649 -26041
rect -741 -26081 -729 -26047
rect -661 -26081 -649 -26047
rect -741 -26087 -649 -26081
rect -463 -26047 -371 -26041
rect -463 -26081 -451 -26047
rect -383 -26081 -371 -26047
rect -463 -26087 -371 -26081
rect -185 -26047 -93 -26041
rect -185 -26081 -173 -26047
rect -105 -26081 -93 -26047
rect -185 -26087 -93 -26081
rect 93 -26047 185 -26041
rect 93 -26081 105 -26047
rect 173 -26081 185 -26047
rect 93 -26087 185 -26081
rect 371 -26047 463 -26041
rect 371 -26081 383 -26047
rect 451 -26081 463 -26047
rect 371 -26087 463 -26081
rect 649 -26047 741 -26041
rect 649 -26081 661 -26047
rect 729 -26081 741 -26047
rect 649 -26087 741 -26081
rect 927 -26047 1019 -26041
rect 927 -26081 939 -26047
rect 1007 -26081 1019 -26047
rect 927 -26087 1019 -26081
rect 1205 -26047 1297 -26041
rect 1205 -26081 1217 -26047
rect 1285 -26081 1297 -26047
rect 1205 -26087 1297 -26081
rect 1483 -26047 1575 -26041
rect 1483 -26081 1495 -26047
rect 1563 -26081 1575 -26047
rect 1483 -26087 1575 -26081
rect 1761 -26047 1853 -26041
rect 1761 -26081 1773 -26047
rect 1841 -26081 1853 -26047
rect 1761 -26087 1853 -26081
rect 2039 -26047 2131 -26041
rect 2039 -26081 2051 -26047
rect 2119 -26081 2131 -26047
rect 2039 -26087 2131 -26081
rect 2317 -26047 2409 -26041
rect 2317 -26081 2329 -26047
rect 2397 -26081 2409 -26047
rect 2317 -26087 2409 -26081
rect 2595 -26047 2687 -26041
rect 2595 -26081 2607 -26047
rect 2675 -26081 2687 -26047
rect 2595 -26087 2687 -26081
<< properties >>
string FIXED_BBOX -2854 -26202 2854 26202
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 260 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
