magic
tech sky130A
timestamp 1697553162
<< end >>
