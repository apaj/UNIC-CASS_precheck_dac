* NGSPICE file created from dac_cell2.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p69_XZX24Q a_n199_n3262# a_n69_n3132# a_n69_2700#
X0 a_n69_2700# a_n69_n3132# a_n199_n3262# sky130_fd_pr__res_xhigh_po_0p69 l=27
C0 a_n69_n3132# a_n199_n3262# 0.805f
C1 a_n69_2700# a_n199_n3262# 0.805f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#1 a_n100_n197# a_100_n100# w_n358_n397#
+ a_n158_n100# VSUBS
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n358_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 w_n358_n397# a_100_n100# 0.1f
C1 w_n358_n397# a_n158_n100# 0.1f
C2 w_n358_n397# a_n100_n197# 0.2f
C3 a_n100_n197# VSUBS 0.282f
C4 w_n358_n397# VSUBS 2.28f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGK6VM a_n100_n297# a_100_n200# w_n358_n497#
+ a_n158_n200# VSUBS
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n358_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
C0 w_n358_n497# a_100_n200# 0.172f
C1 w_n358_n497# a_n158_n200# 0.172f
C2 a_100_n200# a_n158_n200# 0.122f
C3 w_n358_n497# a_n100_n297# 0.2f
C4 a_100_n200# VSUBS 0.105f
C5 a_n158_n200# VSUBS 0.105f
C6 a_n100_n297# VSUBS 0.293f
C7 w_n358_n497# VSUBS 2.81f
.ends

.subckt dac_cell2 vsup vgnd iref vsw iout iout_n vbias
XXR1 vgnd parR sourceM2 sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR2 vgnd parR sourceM2 sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR3 vgnd parR vsup sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR4 vgnd parR vsup sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXM1 iref iref vsup vsup vgnd sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#1
XXM2 iref sourceM3M4 vsup sourceM2 vgnd sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
XXM3 vsw iout vsup sourceM3M4 vgnd sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
XXM4 vbias iout_n vsup sourceM3M4 vgnd sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
C0 vsw vsup 0.161f
C1 iref vsup 1.29f
C2 iout vsw 0.159f
C3 vbias vsup 0.164f
C4 sourceM3M4 vsup 1.61f
C5 sourceM3M4 iout 0.259f
C6 sourceM2 vsup 0.7f
C7 iout vsup 0.233f
C8 iout_n vsup 0.145f
C9 iref sourceM3M4 0.107f
C10 sourceM2 iref 1.36f
C11 iout_n vgnd 0.849f
C12 vbias vgnd 0.528f
C13 iout vgnd 0.379f
C14 sourceM3M4 vgnd 2.06f
C15 vsw vgnd 0.529f
C16 vsup vgnd 15.9f
C17 sourceM2 vgnd 3.21f
C18 iref vgnd 1.63f
C19 parR vgnd 5.35f
.ends

