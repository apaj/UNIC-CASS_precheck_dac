**.subckt tb_esd_cell_tran
x1 net1 pad gate GND esd_cell
V1 net1 GND 3.3
V2 pad GND sine(0 50 1k 0 0 0)
R1 gate GND 100MEG m=1
**** begin user architecture code


.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.param mc_pr_switch=0
*** ANALYSIS TO DO

.tran 10u 5m
.save pad gate

.control
set wr_vecnames
set wr_singlescale

run
******** results filename  ************ nodes to write
wrdata $DEV_PATH/res/tb_esd_cell_tran.res pad gate
.endc


**** end user architecture code
**.ends

* expanding   symbol:  esd_cell.sym # of pins=4
* sym_path: /opt/uniccass/dev/esd_cell/tb/esd_cell.sym
* sch_path: /opt/uniccass/dev/esd_cell/tb/esd_cell.sch
.subckt esd_cell  vsup pad gate vgnd
*.iopin vsup
*.iopin pad
*.iopin vgnd
*.iopin gate
D1 pad vsup sky130_fd_pr__diode_pd2nw_11v0 area=10e+18
D3 gate vsup sky130_fd_pr__diode_pd2nw_05v5 area=0.203e+18
D4 vgnd gate sky130_fd_pr__diode_pw2nd_05v5 area=0.203e+18
XR1 gate pad vgnd sky130_fd_pr__res_high_po W=0.35 L=10 mult=1 m=1
D8 vgnd pad sky130_fd_pr__diode_pw2nd_11v0 area=10e+18
D2 pad vsup sky130_fd_pr__diode_pd2nw_11v0 area=10e+18
D5 pad vsup sky130_fd_pr__diode_pd2nw_11v0 area=10e+18
D6 pad vsup sky130_fd_pr__diode_pd2nw_11v0 area=10e+18
D7 pad vsup sky130_fd_pr__diode_pd2nw_11v0 area=10e+18
D9 vgnd pad sky130_fd_pr__diode_pw2nd_11v0 area=10e+18
D10 vgnd pad sky130_fd_pr__diode_pw2nd_11v0 area=10e+18
D11 vgnd pad sky130_fd_pr__diode_pw2nd_11v0 area=10e+18
D12 vgnd pad sky130_fd_pr__diode_pw2nd_11v0 area=10e+18
.ends

.GLOBAL GND
** flattened .save nodes
.save pad gate
.end
