**.subckt miel21_tb_opamp_op
x1 pow outcm incm incm GND miel21_opamp
V1 incm GND 1.8
V2 pow GND 3.3
R1 outcm GND 1000MEG m=1
**** begin user architecture code


.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.param mc_pr_switch=0
.save incm outcm pow x1.nsources x1.d1 x1.d2 x1.bias
.save @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[id]
.save @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[id]
.save @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[id]
.save @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[id]
.save @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[id]
.save @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[id]
.save @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[id]
.save @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[id] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[gm] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[gm] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[gm] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vdsat] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vdsat] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vdsat] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vds] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vds] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vds] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vgs] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vgs] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vgs] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vth] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vth] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vth]
.op

.control
set wr_vecnames
set wr_singlescale

run

wrdata miel21_tb_opamp_op.res incm outcm pow x1.nsources x1.d1 x1.d2 x1.bias
+ @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[id] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[id] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[id]
+ @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[id] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[id] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[id]
+ @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[id] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[id] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[gm]
+ @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[gm]
+ @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[gm] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[gm]
+ @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[gm] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
+ @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
+ @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vdsat] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vdsat] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
+ @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vds]
+ @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vds]
+ @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vds] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vds] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs]
+ @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vgs]
+ @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vgs] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vgs]
+ @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vgs] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vth]
+ @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vth]
+ @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vth] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vth] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vth]
.endc


**** end user architecture code
**.ends

* expanding   symbol:  miel21_opamp.sym # of pins=5
* sym_path: /opt/uniccass/dev/opamp/miel21_opamp.sym
* sch_path: /opt/uniccass/dev/opamp/miel21_opamp.sch
.subckt miel21_opamp  power outSingle inPos inNeg ground
*.ipin inPos
*.ipin inNeg
*.opin outSingle
*.iopin power
*.iopin ground
XM6 d1 d1 power power sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=21 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 d2 d1 power power sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=21 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 outSingle d2 power power sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=260 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM1 d1 inPos nsources ground sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM2 d2 inNeg nsources ground sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 bias bias ground ground sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 nsources bias ground ground sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM5 outSingle bias ground ground sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=48 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XR1 bias net2 ground sky130_fd_pr__res_xhigh_po_0p69 L=6 mult=1 m=1
XC1 outSingle d2 sky130_fd_pr__cap_mim_m3_1 W=10 L=14 MF=1 m=1
XR2 net2 net1 ground sky130_fd_pr__res_xhigh_po_0p69 L=6 mult=1 m=1
XR3 net1 power ground sky130_fd_pr__res_xhigh_po_0p69 L=6 mult=1 m=1
.ends

.GLOBAL GND
** flattened .save nodes
.save incm outcm pow x1.nsources x1.d1 x1.d2 x1.bias
.save @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[id]
.save @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[id]
.save @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[id]
.save @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[id]
.save @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[id]
.save @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[id]
.save @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[id]
.save @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[id] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[gm] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[gm] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[gm] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[gm] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vdsat] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vdsat] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vdsat] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vdsat] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vds] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vds] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vds] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vds] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vgs] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vgs] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vgs] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vgs] @m.x1.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm2.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm3.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm4.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm5.msky130_fd_pr__nfet_g5v0d10v5[vth] @m.x1.xm6.msky130_fd_pr__pfet_g5v0d10v5[vth] @m.x1.xm7.msky130_fd_pr__pfet_g5v0d10v5[vth] @m.x1.xm8.msky130_fd_pr__pfet_g5v0d10v5[vth]
.end
