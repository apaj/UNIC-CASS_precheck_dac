magic
tech sky130A
magscale 1 2
timestamp 1698257525
<< psubdiff >>
rect 7180 7410 8510 7490
rect 7180 6550 7280 7410
rect 8460 6550 8510 7410
rect 7180 6480 8510 6550
<< psubdiffcont >>
rect 7280 6550 8460 7410
<< viali >>
rect 7170 7410 8510 7500
rect 7170 6550 7280 7410
rect 7280 6550 8460 7410
rect 8460 6550 8510 7410
rect 15306 6596 15352 6754
rect 7170 6480 8510 6550
rect 15314 6172 15360 6330
rect 15330 5740 15376 5898
rect 15314 5318 15360 5476
rect -194 -5092 18 -4882
rect 8062 -9386 8104 -8742
rect 8056 -10280 8098 -9636
rect 8046 -11180 8088 -10536
rect -6552 -12600 -5916 -11902
rect 8046 -12078 8088 -11434
rect -10190 -14018 -10144 -12798
rect -10198 -15476 -10160 -14258
rect -10204 -16964 -10166 -15746
rect -10230 -18428 -10192 -17210
<< metal1 >>
rect -10402 11398 -4450 11412
rect -10402 11352 -4446 11398
rect -23348 11114 -21974 11246
rect -23348 9058 -22894 11114
rect -22328 9058 -21974 11114
rect -10402 10768 -10362 11352
rect -9028 10768 -4446 11352
rect -10402 10726 -4446 10768
rect -10402 10718 -4450 10726
rect -16192 9606 -14820 9726
rect 9676 9638 10016 11634
rect -16192 9124 -16040 9606
rect -23348 5308 -21974 9058
rect -16262 8992 -16040 9124
rect -14996 8992 -14820 9606
rect 5352 9630 10016 9638
rect 5352 9190 5356 9630
rect 6124 9190 10016 9630
rect 5352 9172 10016 9190
rect -16262 8972 -16030 8992
rect -15892 8972 -14820 8992
rect -16262 8960 -14820 8972
rect -16262 8954 -15840 8960
rect -21780 8772 -21496 8838
rect -21780 8552 -21746 8772
rect -21538 8552 -21496 8772
rect -21780 8500 -21496 8552
rect -2746 8542 -2286 8566
rect -8024 8480 -7090 8482
rect -2746 8480 -2728 8542
rect -8024 8462 -2728 8480
rect -8024 8046 -7980 8462
rect -7220 8046 -2728 8462
rect -8024 8028 -2728 8046
rect -2310 8028 -2286 8542
rect -8024 8018 -2286 8028
rect -7180 8012 -2286 8018
rect -2746 8010 -2286 8012
rect 9440 7580 10002 9172
rect 7060 7500 10002 7580
rect -3386 7294 -1396 7370
rect -3386 6950 -3284 7294
rect -2872 6950 -1396 7294
rect -3386 6896 -1396 6950
rect -1240 7200 -644 7232
rect -1240 6918 -1206 7200
rect -670 6918 -644 7200
rect -1596 6886 -1406 6896
rect -1240 6892 -644 6918
rect -494 6596 -286 7462
rect 3796 7316 4888 7322
rect -34 6996 4888 7316
rect -6682 6594 -6638 6596
rect -5800 6594 -286 6596
rect -6682 6576 -286 6594
rect -6682 6318 -6654 6576
rect -5824 6318 -286 6576
rect -6682 6298 -286 6318
rect -23348 3314 -23060 5308
rect -22202 3314 -21974 5308
rect 2774 5946 3260 5972
rect 2774 5542 2804 5946
rect 3238 5542 3260 5946
rect -10402 4990 -4374 5080
rect -10402 4406 -10368 4990
rect -9034 4406 -4374 4990
rect -10402 4344 -4374 4406
rect -16122 3808 -14932 3856
rect -16122 3472 -15896 3808
rect -16168 3362 -15896 3472
rect -23348 -308 -21974 3314
rect -16176 3188 -15896 3362
rect -14952 3188 -14932 3808
rect -16176 3182 -14932 3188
rect -16168 3178 -14932 3182
rect -16168 3176 -15624 3178
rect -21820 3012 -21436 3064
rect -21820 2750 -21738 3012
rect -21498 2750 -21436 3012
rect -21820 2682 -21436 2750
rect 2774 2172 3260 5542
rect -8028 1672 -4638 1674
rect -8028 1614 -4240 1672
rect -8028 1106 -8000 1614
rect -7240 1106 -4240 1614
rect -8028 1046 -4240 1106
rect -7180 1042 -4240 1046
rect 3796 292 4888 6996
rect 7060 6480 7170 7500
rect 8510 6824 10002 7500
rect 8510 6754 15378 6824
rect 8510 6596 15306 6754
rect 15352 6596 15378 6754
rect 16702 6756 21528 6758
rect 8510 6480 15378 6596
rect 7060 6372 15378 6480
rect 7060 6370 9520 6372
rect 15284 6330 15378 6372
rect 15284 6172 15314 6330
rect 15360 6172 15378 6330
rect 15284 5908 15378 6172
rect 15284 5898 15390 5908
rect 15284 5740 15330 5898
rect 15376 5740 15390 5898
rect 15284 5732 15390 5740
rect 15284 5476 15378 5732
rect 15284 5318 15314 5476
rect 15360 5318 15378 5476
rect 15440 5366 15882 6724
rect 16702 6212 22178 6756
rect 16722 5848 17182 5852
rect 16720 5358 17182 5848
rect 15284 5280 15378 5318
rect 16722 4972 17182 5358
rect -2306 172 -1712 200
rect -23348 -2302 -23146 -308
rect -22288 -2302 -21974 -308
rect -4432 38 -2442 142
rect -4432 -192 -4270 38
rect -3964 -192 -2442 38
rect -2306 -126 -2276 172
rect -1742 -126 -1712 172
rect -2306 -146 -1712 -126
rect -4432 -332 -2442 -192
rect -6684 -432 -5734 -428
rect -1464 -432 -1256 258
rect -734 -28 4888 292
rect -6684 -468 -1256 -432
rect -6684 -918 -6654 -468
rect -5826 -918 -1256 -468
rect -6684 -948 -1256 -918
rect -6684 -950 -5734 -948
rect 2756 -1054 3154 -1030
rect 2756 -1452 2784 -1054
rect 3130 -1452 3154 -1054
rect -10402 -1602 -2286 -1546
rect -10402 -2186 -10364 -1602
rect -9030 -2186 -2286 -1602
rect -10402 -2236 -2286 -2186
rect -16100 -2278 -15638 -2268
rect -23348 -5978 -21974 -2302
rect -16240 -2458 -15638 -2278
rect -21844 -2644 -21430 -2582
rect -21844 -2992 -21776 -2644
rect -21474 -2992 -21430 -2644
rect -21844 -3104 -21430 -2992
rect -23348 -7972 -23146 -5978
rect -22288 -7972 -21974 -5978
rect -16100 -5116 -15638 -2458
rect 2756 -3898 3154 -1452
rect -8026 -4898 -2330 -4880
rect -252 -4882 62 -4854
rect -8026 -4900 -2328 -4898
rect -16100 -5210 -12432 -5116
rect -8026 -5162 -8014 -4900
rect -7196 -4920 -2328 -4900
rect -7196 -5142 -3234 -4920
rect -2350 -5142 -2328 -4920
rect -7196 -5154 -2328 -5142
rect -252 -5092 -194 -4882
rect 18 -5092 62 -4882
rect -7196 -5162 -2330 -5154
rect -8026 -5176 -2330 -5162
rect -7180 -5178 -2330 -5176
rect -252 -5186 62 -5092
rect -16100 -6182 -14338 -5210
rect -16116 -6634 -14338 -6182
rect -16100 -6644 -14338 -6634
rect -16096 -6672 -14338 -6644
rect -12486 -6672 -12432 -5210
rect -16096 -6746 -12432 -6672
rect -23348 -11648 -21974 -7972
rect -16130 -7294 -14224 -7158
rect -16130 -7978 -15680 -7294
rect -16204 -8150 -15680 -7978
rect -21830 -8314 -21448 -8276
rect -21830 -8656 -21796 -8314
rect -21484 -8656 -21448 -8314
rect -16130 -8362 -15680 -8150
rect -14350 -8362 -14224 -7294
rect -1198 -7484 792 -7446
rect -1198 -7842 -1100 -7484
rect -672 -7842 792 -7484
rect -1198 -7920 792 -7842
rect 1010 -7520 1030 -7500
rect 1010 -7540 1604 -7520
rect 1010 -7852 1026 -7540
rect 1578 -7852 1604 -7540
rect 1010 -7872 1604 -7852
rect -16130 -8462 -14224 -8362
rect -6678 -8056 -5694 -8050
rect -6678 -8060 -5252 -8056
rect -6678 -8062 -3794 -8060
rect 1770 -8062 1978 -7234
rect 3796 -7458 4888 -28
rect 6706 4460 17182 4972
rect 6706 -1082 7894 4460
rect 16722 4458 17182 4460
rect 21542 2346 22178 6212
rect 21542 2256 22744 2346
rect 21542 296 21716 2256
rect 22146 716 22744 2256
rect 21538 260 21716 296
rect 22158 296 22744 716
rect 22158 262 22746 296
rect 22146 260 22746 262
rect 21538 -824 22746 260
rect 6706 -1744 9874 -1082
rect 2174 -7778 4888 -7458
rect -6678 -8072 1978 -8062
rect -6678 -8546 -6662 -8072
rect -5828 -8546 1978 -8072
rect -6678 -8570 1978 -8546
rect -6674 -8574 1978 -8570
rect -5800 -8578 1978 -8574
rect 2240 -8404 2742 -8384
rect -5274 -8586 -3794 -8578
rect -21830 -8706 -21448 -8656
rect 2240 -8812 2266 -8404
rect 2720 -8812 2742 -8404
rect -10402 -9330 -1072 -9316
rect -10402 -9374 -1070 -9330
rect -10402 -9958 -10356 -9374
rect -9022 -9958 -1070 -9374
rect -10402 -10002 -1070 -9958
rect -10402 -10006 -1072 -10002
rect -23348 -13366 -23050 -11648
rect -23392 -13642 -23050 -13366
rect -22192 -13642 -21974 -11648
rect 632 -11522 988 -11498
rect 632 -11706 664 -11522
rect 958 -11706 988 -11522
rect 2240 -11684 2742 -8812
rect 632 -11736 988 -11706
rect -16146 -11792 -15592 -11788
rect -16146 -11884 -5826 -11792
rect -16146 -12630 -6584 -11884
rect -5912 -12630 -5826 -11884
rect -16146 -12686 -5826 -12630
rect -16146 -13332 -15592 -12686
rect -10250 -12798 -10126 -12782
rect -16146 -13588 -15590 -13332
rect -23392 -13766 -21974 -13642
rect -16158 -13760 -15590 -13588
rect -23392 -18660 -22034 -13766
rect -21868 -13936 -21464 -13886
rect -21868 -14312 -21810 -13936
rect -21530 -14312 -21464 -13936
rect -21868 -14370 -21464 -14312
rect -10250 -14018 -10190 -12798
rect -10144 -14018 -10126 -12798
rect -10250 -14048 -10126 -14018
rect -10250 -14258 -10128 -14048
rect -10250 -15476 -10198 -14258
rect -10160 -15476 -10128 -14258
rect -10250 -15746 -10128 -15476
rect -10250 -16964 -10204 -15746
rect -10166 -16964 -10128 -15746
rect -10250 -17210 -10128 -16964
rect -10250 -18426 -10230 -17210
rect -10252 -18428 -10230 -18426
rect -10192 -18428 -10128 -17210
rect -10096 -18392 -9626 -12816
rect -9382 -12936 -7184 -12816
rect -9382 -14352 -7988 -12936
rect -7260 -14352 -7184 -12936
rect -9382 -14482 -7184 -14352
rect -9370 -15424 -8944 -14482
rect -7218 -14484 -7184 -14482
rect -9404 -17982 -8978 -15788
rect 3796 -16014 4888 -7778
rect 6718 -1756 9874 -1744
rect 6718 -1758 8336 -1756
rect 6718 -7718 7542 -1758
rect 8656 -4340 10006 -2124
rect 8656 -5132 8818 -4340
rect 9770 -5132 10006 -4340
rect 8656 -6082 10006 -5132
rect 6718 -8384 9316 -7718
rect 6718 -8386 8218 -8384
rect 8012 -8716 8104 -8646
rect 8012 -8742 8114 -8716
rect 8012 -9386 8062 -8742
rect 8104 -9386 8114 -8742
rect 8012 -9404 8114 -9386
rect 8012 -9636 8104 -9404
rect 8012 -10254 8056 -9636
rect 5364 -10280 8056 -10254
rect 8098 -10280 8104 -9636
rect 5364 -10292 8104 -10280
rect 5364 -10740 5390 -10292
rect 6124 -10536 8104 -10292
rect 6124 -10740 8046 -10536
rect 5364 -10772 8046 -10740
rect 8012 -11180 8046 -10772
rect 8088 -11180 8104 -10536
rect 8012 -11434 8104 -11180
rect 8012 -12078 8046 -11434
rect 8088 -12078 8104 -11434
rect 8170 -12070 8622 -8776
rect 8876 -10266 9316 -8384
rect 8012 -12136 8104 -12078
rect 8858 -12234 9298 -10580
rect 25476 -11374 26284 -11248
rect 14806 -11578 15404 -11504
rect 25476 -11506 25590 -11374
rect 14806 -11942 14848 -11578
rect 15332 -11942 15404 -11578
rect 14806 -12034 15404 -11942
rect 21154 -11948 25590 -11506
rect 8810 -16010 9304 -12234
rect 14806 -12278 15766 -12034
rect 25476 -12060 25590 -11948
rect 26142 -12060 26284 -11374
rect 25476 -12172 26284 -12060
rect 14806 -12280 15404 -12278
rect 7512 -16014 9304 -16010
rect 1536 -16702 2132 -16688
rect -650 -16822 1340 -16794
rect -650 -17204 -582 -16822
rect -126 -17204 1340 -16822
rect 1536 -17032 1550 -16702
rect 2114 -17032 2132 -16702
rect 1536 -17038 2132 -17032
rect -650 -17268 1340 -17204
rect -6678 -17396 -4624 -17392
rect -6678 -17408 -4618 -17396
rect 2372 -17408 2580 -16522
rect 3796 -16686 9304 -16014
rect 2762 -16986 9304 -16686
rect 2762 -17006 4888 -16986
rect 7512 -16990 9304 -16986
rect 7512 -16994 9286 -16990
rect -6678 -17424 2580 -17408
rect -6678 -17900 -6640 -17424
rect -5834 -17900 2580 -17424
rect -6678 -17924 2580 -17900
rect -6678 -17930 -4618 -17924
rect -6678 -17932 -5796 -17930
rect -9420 -18344 -8974 -17982
rect -10252 -18654 -10128 -18428
rect -9420 -18540 -7508 -18344
rect -9420 -18654 -9252 -18540
rect -10254 -18660 -9252 -18654
rect -23392 -19020 -9252 -18660
rect -7716 -19020 -7508 -18540
rect -23392 -19162 -7508 -19020
rect -21944 -19170 -7520 -19162
rect -10254 -19172 -7520 -19170
<< via1 >>
rect -22894 9058 -22328 11114
rect -10362 10768 -9028 11352
rect -16040 8992 -14996 9606
rect 5356 9190 6124 9630
rect -16030 8972 -15892 8992
rect -21746 8552 -21538 8772
rect -7980 8046 -7220 8462
rect -2728 8028 -2310 8542
rect -3284 6950 -2872 7294
rect -1206 6918 -670 7200
rect -6654 6318 -5824 6576
rect -23060 3314 -22202 5308
rect 2804 5542 3238 5946
rect -10368 4406 -9034 4990
rect -15896 3188 -14952 3808
rect -21738 2750 -21498 3012
rect -8000 1106 -7240 1614
rect -23146 -2302 -22288 -308
rect -4270 -192 -3964 38
rect -2276 -126 -1742 172
rect -6654 -918 -5826 -468
rect 2784 -1452 3130 -1054
rect -10364 -2186 -9030 -1602
rect -21776 -2992 -21474 -2644
rect -23146 -7972 -22288 -5978
rect -8014 -5162 -7196 -4900
rect -3234 -5142 -2350 -4920
rect -194 -5092 18 -4882
rect -14338 -6672 -12486 -5210
rect -21796 -8656 -21484 -8314
rect -15680 -8362 -14350 -7294
rect -1100 -7842 -672 -7484
rect 1026 -7852 1578 -7540
rect 21716 716 22146 2256
rect 21716 262 22158 716
rect 21716 260 22146 262
rect -6662 -8546 -5828 -8072
rect 2266 -8812 2720 -8404
rect -10356 -9958 -9022 -9374
rect -23050 -13642 -22192 -11648
rect 664 -11706 958 -11522
rect -6584 -11902 -5912 -11884
rect -6584 -12600 -6552 -11902
rect -6552 -12600 -5916 -11902
rect -5916 -12600 -5912 -11902
rect -6584 -12630 -5912 -12600
rect -21810 -14312 -21530 -13936
rect -7988 -14352 -7260 -12936
rect 8818 -5132 9770 -4340
rect 5390 -10740 6124 -10292
rect 14848 -11942 15332 -11578
rect 25590 -12060 26142 -11374
rect -582 -17204 -126 -16822
rect 1550 -17032 2114 -16702
rect -6640 -17900 -5834 -17424
rect -9252 -19020 -7716 -18540
<< metal2 >>
rect 13742 14424 24242 14434
rect -10406 14418 24242 14424
rect -26762 14064 24242 14418
rect -26762 13028 -5488 14064
rect -4428 13028 24242 14064
rect -26762 12854 24242 13028
rect -26762 12298 -9024 12854
rect -26732 8248 -24706 12298
rect -10406 11420 -9024 12298
rect 13268 12756 24242 12854
rect -10406 11352 -8978 11420
rect -23088 11218 -22176 11230
rect -23088 11114 -21330 11218
rect -23088 9058 -22894 11114
rect -22328 9058 -21330 11114
rect -10406 10768 -10362 11352
rect -9028 10768 -8978 11352
rect -10406 10714 -8978 10768
rect -23088 8932 -21330 9058
rect -16128 9606 -14916 9638
rect -16128 8992 -16040 9606
rect -14996 8992 -14916 9606
rect -10402 9220 -8978 10714
rect 5352 9630 6142 9640
rect -10402 9036 -8976 9220
rect -16128 8968 -16036 8992
rect -15860 8968 -14916 8992
rect -16128 8960 -14916 8968
rect -16052 8956 -15840 8960
rect -23088 8918 -22176 8932
rect -21770 8776 -21512 8806
rect -21770 8546 -21752 8776
rect -21534 8546 -21512 8776
rect -21770 8512 -21512 8546
rect -26732 5940 -21492 8248
rect -10398 6528 -8976 9036
rect 5352 9190 5356 9630
rect 6124 9190 6142 9630
rect -2746 8542 -2286 8566
rect -10402 6488 -8976 6528
rect -8026 8462 -7180 8480
rect -8026 8046 -7980 8462
rect -7220 8046 -7180 8462
rect -26732 2532 -24706 5940
rect -23210 5308 -21346 5458
rect -23210 3314 -23060 5308
rect -22202 3314 -21346 5308
rect -10402 4990 -8978 6488
rect -10402 4406 -10368 4990
rect -9034 4406 -8978 4990
rect -23210 3218 -21346 3314
rect -22942 3176 -21346 3218
rect -15936 3808 -14940 3828
rect -15936 3188 -15896 3808
rect -14952 3188 -14940 3808
rect -15896 3180 -15630 3188
rect -21786 3032 -21470 3046
rect -21786 2724 -21774 3032
rect -21482 2724 -21470 3032
rect -21786 2716 -21470 2724
rect -26732 224 -21424 2532
rect -26732 -3148 -24706 224
rect -23318 -308 -21454 -222
rect -23318 -2302 -23146 -308
rect -22288 -2302 -21454 -308
rect -23318 -2462 -21454 -2302
rect -10402 -1602 -8978 4406
rect -10402 -2186 -10364 -1602
rect -9030 -2186 -8978 -1602
rect -21844 -2630 -21432 -2580
rect -21844 -2998 -21800 -2630
rect -21464 -2998 -21432 -2630
rect -21844 -3042 -21432 -2998
rect -26732 -5456 -21402 -3148
rect -14406 -5210 -12466 -5166
rect -26732 -8842 -24706 -5456
rect -23306 -5978 -21442 -5894
rect -23306 -7972 -23146 -5978
rect -22288 -7972 -21442 -5978
rect -14406 -6672 -14338 -5210
rect -12486 -6672 -12466 -5210
rect -14406 -6698 -12466 -6672
rect -23306 -8134 -21442 -7972
rect -15698 -7294 -14270 -7240
rect -21826 -8298 -21446 -8274
rect -21826 -8658 -21810 -8298
rect -21472 -8658 -21446 -8298
rect -15698 -8362 -15680 -7294
rect -14350 -8362 -14270 -7294
rect -15698 -8426 -14270 -8362
rect -21826 -8678 -21446 -8658
rect -26732 -11150 -21436 -8842
rect -10402 -9374 -8978 -2186
rect -10402 -9958 -10356 -9374
rect -9022 -9958 -8978 -9374
rect -10402 -10010 -8978 -9958
rect -8026 1614 -7180 8046
rect -2746 8028 -2728 8542
rect -2310 8028 -2286 8542
rect -2746 8010 -2286 8028
rect -3752 7294 -2706 7372
rect -3752 7290 -3284 7294
rect -3752 6948 -3710 7290
rect -3370 6950 -3284 7290
rect -2872 6950 -2706 7294
rect -3370 6948 -2706 6950
rect -3752 6890 -2706 6948
rect -1240 7200 -644 7232
rect -1240 6918 -1206 7200
rect -670 6918 -644 7200
rect -1240 6892 -644 6918
rect -6678 6576 -5800 6596
rect -6678 6318 -6654 6576
rect -5824 6318 -5800 6576
rect -6678 1730 -5800 6318
rect -1064 5972 -644 6892
rect 5352 5972 6142 9190
rect -1074 5968 6142 5972
rect -1074 5946 6148 5968
rect -1074 5542 2804 5946
rect 3238 5542 6148 5946
rect -1074 5504 6148 5542
rect -1064 5496 -644 5504
rect -6684 1654 -5798 1730
rect -8026 1106 -8000 1614
rect -7240 1106 -7180 1614
rect -8026 -4900 -7180 1106
rect -8026 -5162 -8014 -4900
rect -7196 -5162 -7180 -4900
rect -8026 -10388 -7180 -5162
rect -6678 -468 -5800 1654
rect -4628 1062 -4150 1672
rect -2306 172 -1712 200
rect -4674 56 -3788 148
rect -4674 -308 -4620 56
rect -4258 38 -3788 56
rect -3964 -192 -3788 38
rect -2306 -126 -2276 172
rect -1742 -126 -1712 172
rect -2306 -146 -1712 -126
rect -4258 -308 -3788 -192
rect -4674 -326 -3788 -308
rect -6678 -918 -6654 -468
rect -5826 -918 -5800 -468
rect -6678 -2268 -5800 -918
rect -2132 -1026 -1712 -146
rect 5362 -1026 6148 5504
rect 13268 4164 14040 12756
rect 10556 3264 14044 4164
rect 21648 2336 22738 2346
rect 21538 2256 22738 2336
rect 21538 260 21716 2256
rect 22146 716 22196 2256
rect 22158 714 22196 716
rect 22626 828 22738 2256
rect 22158 262 22194 714
rect 22146 260 22194 262
rect 22626 296 22742 828
rect 22626 260 22746 296
rect 21538 258 22194 260
rect 22622 258 22746 260
rect 21538 -824 22746 258
rect -2150 -1054 6148 -1026
rect -2150 -1452 2784 -1054
rect 3130 -1452 6148 -1054
rect -2150 -1494 6148 -1452
rect -2132 -1502 -1712 -1494
rect -6678 -4836 -5812 -2268
rect 5362 -3364 6148 -1494
rect 7168 -3364 8644 -3360
rect 5362 -3964 11088 -3364
rect 5362 -3972 7542 -3964
rect 8288 -3972 11088 -3964
rect -6678 -8072 -5800 -4836
rect -254 -4882 66 -4852
rect -254 -4898 -194 -4882
rect -3248 -4920 -194 -4898
rect -3248 -5142 -3234 -4920
rect -2350 -5092 -194 -4920
rect 18 -5092 66 -4882
rect -2350 -5142 66 -5092
rect -3248 -5154 66 -5142
rect -2566 -5158 66 -5154
rect -254 -5188 66 -5158
rect -1388 -7484 -652 -7444
rect -1388 -7502 -1100 -7484
rect -1388 -7894 -1298 -7502
rect -672 -7842 -652 -7484
rect 1178 -7520 1610 -7514
rect -868 -7894 -652 -7842
rect 1010 -7540 1610 -7520
rect 1010 -7852 1026 -7540
rect 1578 -7852 1610 -7540
rect 1010 -7872 1610 -7852
rect -1388 -7932 -652 -7894
rect -6678 -8546 -6662 -8072
rect -5828 -8546 -5800 -8072
rect -8026 -10678 -7182 -10388
rect -6678 -10418 -5800 -8546
rect 1124 -8382 1610 -7872
rect 5362 -8382 6148 -3972
rect 10498 -4102 11088 -3972
rect 8656 -4340 10002 -4124
rect 8656 -5132 8818 -4340
rect 9770 -5132 10002 -4340
rect 8656 -5206 10002 -5132
rect 8656 -6010 8818 -5206
rect 9778 -6010 10002 -5206
rect 8656 -6082 10002 -6010
rect 1124 -8404 6148 -8382
rect 1124 -8812 2266 -8404
rect 2720 -8812 6148 -8404
rect 1124 -8850 6148 -8812
rect 1124 -8856 1610 -8850
rect 1124 -8860 1592 -8856
rect -26732 -14450 -24706 -11150
rect -8026 -11280 -7180 -10678
rect -23220 -11648 -21356 -11500
rect -23220 -13642 -23050 -11648
rect -22192 -13642 -21356 -11648
rect -23220 -13740 -21356 -13642
rect -8048 -11512 -7180 -11280
rect -6680 -11380 -5800 -10418
rect -8048 -11720 -8016 -11512
rect -7190 -11720 -7180 -11512
rect -8048 -12936 -7180 -11720
rect -21844 -13928 -21498 -13910
rect -21844 -14312 -21824 -13928
rect -21524 -14312 -21498 -13928
rect -21844 -14338 -21498 -14312
rect -8048 -14352 -7988 -12936
rect -7260 -14352 -7180 -12936
rect -26732 -14472 -21612 -14450
rect -26732 -16696 -21354 -14472
rect -8048 -14482 -7180 -14352
rect -6678 -11884 -5800 -11380
rect 5362 -10292 6148 -8850
rect 23308 -9074 24228 12756
rect 5362 -10740 5390 -10292
rect 6124 -10740 6148 -10292
rect 626 -11518 980 -11498
rect 626 -11706 656 -11518
rect 960 -11706 980 -11518
rect 626 -11730 980 -11706
rect -6678 -12630 -6584 -11884
rect -5912 -12630 -5800 -11884
rect -25304 -16762 -21354 -16696
rect -25304 -16774 -21612 -16762
rect -6678 -17424 -5800 -12630
rect 1536 -16702 2132 -16688
rect -1118 -16744 -502 -16734
rect -1118 -16808 -72 -16744
rect -1118 -17200 -1018 -16808
rect -574 -16822 -72 -16808
rect -1118 -17204 -582 -17200
rect -126 -17204 -72 -16822
rect 1536 -17032 1550 -16702
rect 2114 -17032 2132 -16702
rect 1536 -17038 2132 -17032
rect -1118 -17276 -72 -17204
rect -688 -17286 -72 -17276
rect -6678 -17900 -6640 -17424
rect -5834 -17900 -5800 -17424
rect -6678 -17932 -5800 -17900
rect 1698 -17904 2130 -17038
rect 5362 -17870 6148 -10740
rect 20928 -11296 24228 -9074
rect 25528 -11300 26264 -11264
rect 14838 -11572 15344 -11558
rect 14838 -11948 14846 -11572
rect 15334 -11948 15344 -11572
rect 14838 -11964 15344 -11948
rect 20996 -14374 24222 -12000
rect 25528 -12096 25552 -11300
rect 26182 -12096 26264 -11300
rect 25528 -12156 26264 -12096
rect 23260 -17870 24216 -14374
rect 5358 -17904 24216 -17870
rect 1688 -18350 24216 -17904
rect -9428 -18522 24216 -18350
rect -9428 -18540 -6384 -18522
rect -9428 -19020 -9252 -18540
rect -7716 -19020 -6384 -18540
rect -9428 -19054 -6384 -19020
rect -5662 -19054 24216 -18522
rect -9428 -19146 24216 -19054
rect -9428 -19150 23940 -19146
rect 6030 -19156 6146 -19150
<< via2 >>
rect -5488 13028 -4428 14064
rect -16040 8992 -14996 9606
rect -16036 8972 -16030 8992
rect -16030 8972 -15892 8992
rect -15892 8972 -15860 8992
rect -16036 8968 -15860 8972
rect -21752 8772 -21534 8776
rect -21752 8552 -21746 8772
rect -21746 8552 -21538 8772
rect -21538 8552 -21534 8772
rect -21752 8546 -21534 8552
rect -15896 3188 -14952 3808
rect -21774 3012 -21482 3032
rect -21774 2750 -21738 3012
rect -21738 2750 -21498 3012
rect -21498 2750 -21482 3012
rect -21774 2724 -21482 2750
rect -21800 -2644 -21464 -2630
rect -21800 -2992 -21776 -2644
rect -21776 -2992 -21474 -2644
rect -21474 -2992 -21464 -2644
rect -21800 -2998 -21464 -2992
rect -14338 -6672 -12486 -5210
rect -21810 -8314 -21472 -8298
rect -21810 -8656 -21796 -8314
rect -21796 -8656 -21484 -8314
rect -21484 -8656 -21472 -8314
rect -21810 -8658 -21472 -8656
rect -15680 -8362 -14350 -7294
rect -3710 6948 -3370 7290
rect -4620 38 -4258 56
rect -4620 -192 -4270 38
rect -4270 -192 -4258 38
rect -4620 -308 -4258 -192
rect 22196 714 22626 2256
rect 22194 260 22626 714
rect 22194 258 22622 260
rect -1298 -7842 -1100 -7502
rect -1100 -7842 -868 -7502
rect -1298 -7894 -868 -7842
rect 8818 -6010 9778 -5206
rect -8016 -11720 -7190 -11512
rect -21824 -13936 -21524 -13928
rect -21824 -14312 -21810 -13936
rect -21810 -14312 -21530 -13936
rect -21530 -14312 -21524 -13936
rect 656 -11522 960 -11518
rect 656 -11706 664 -11522
rect 664 -11706 958 -11522
rect 958 -11706 960 -11522
rect -1018 -16822 -574 -16808
rect -1018 -17200 -582 -16822
rect -582 -17200 -574 -16822
rect 14846 -11578 15334 -11572
rect 14846 -11942 14848 -11578
rect 14848 -11942 15332 -11578
rect 15332 -11942 15334 -11578
rect 14846 -11948 15334 -11942
rect 25552 -11374 26182 -11300
rect 25552 -12060 25590 -11374
rect 25590 -12060 26142 -11374
rect 26142 -12060 26182 -11374
rect 25552 -12096 26182 -12060
rect -6384 -19054 -5662 -18522
<< metal3 >>
rect -5830 14064 -4152 18344
rect -5830 13028 -5488 14064
rect -4428 13028 -4152 14064
rect -5830 12834 -4152 13028
rect -16088 9606 -14772 9870
rect -16088 8992 -16040 9606
rect -14996 8992 -14772 9606
rect -16088 8968 -16036 8992
rect -15860 8968 -14772 8992
rect -27912 8932 -21954 8958
rect -27912 8776 -21408 8932
rect -27912 8546 -21752 8776
rect -21534 8546 -21408 8776
rect -27912 8346 -21408 8546
rect -27366 8320 -21408 8346
rect -16088 7670 -14772 8968
rect -16088 7290 -2720 7670
rect -16088 6948 -3710 7290
rect -3370 6948 -2720 7290
rect -16088 6776 -2720 6948
rect -15908 3808 -14916 3916
rect -28028 3032 -21434 3192
rect -15908 3188 -15896 3808
rect -14952 3478 -14916 3808
rect -14952 3188 -14908 3478
rect -15908 3086 -14908 3188
rect -28028 2724 -21774 3032
rect -21482 2724 -21434 3032
rect -28028 2436 -21434 2724
rect -15904 380 -14908 3086
rect 22024 2256 25932 2500
rect 22024 714 22196 2256
rect -15904 378 -14060 380
rect -15904 370 -4258 378
rect -15904 56 -3706 370
rect -15904 -308 -4620 56
rect -4258 -308 -3706 56
rect -15904 -396 -3706 -308
rect -15892 -398 -3706 -396
rect -15892 -400 -14060 -398
rect -11910 -408 -3706 -398
rect 22024 258 22194 714
rect 22626 260 25932 2256
rect 22622 258 25932 260
rect -11910 -410 -3794 -408
rect 22024 -1160 25932 258
rect -27890 -2630 -21420 -2524
rect -27890 -2998 -21800 -2630
rect -21464 -2998 -21420 -2630
rect -27890 -3416 -21420 -2998
rect -14388 -5210 -12412 -5030
rect -14388 -6672 -14338 -5210
rect -12486 -6672 -12412 -5210
rect 8610 -5206 15540 -4988
rect 8610 -6010 8818 -5206
rect 9778 -6010 15540 -5206
rect 8610 -6604 15540 -6010
rect -14388 -6762 -12412 -6672
rect -15716 -7294 -14172 -7114
rect -27744 -8298 -21418 -8132
rect -27744 -8658 -21810 -8298
rect -21472 -8658 -21418 -8298
rect -15716 -8362 -15680 -7294
rect -14350 -8362 -14172 -7294
rect -13676 -7262 -12412 -6762
rect 14798 -6622 15540 -6604
rect -13676 -7264 -868 -7262
rect -13676 -7502 -534 -7264
rect -13676 -7894 -1298 -7502
rect -868 -7894 -534 -7502
rect -13676 -8100 -534 -7894
rect -888 -8102 -534 -8100
rect -15716 -8444 -14172 -8362
rect -27744 -8934 -21418 -8658
rect -15744 -8464 -11260 -8444
rect -15744 -9952 -11132 -8464
rect -22160 -13928 -21432 -13848
rect -22160 -14312 -21824 -13928
rect -21524 -14312 -21432 -13928
rect -22160 -19764 -21432 -14312
rect -13502 -16188 -11132 -9952
rect -8026 -11512 984 -11500
rect -8026 -11720 -8016 -11512
rect -7190 -11518 984 -11512
rect -7190 -11706 656 -11518
rect 960 -11706 984 -11518
rect -7190 -11720 984 -11706
rect -8026 -11726 984 -11720
rect -8026 -11728 -7180 -11726
rect -2734 -11730 984 -11726
rect 14798 -11572 15542 -6622
rect 14798 -11948 14846 -11572
rect 15334 -11948 15542 -11572
rect 14798 -11970 15542 -11948
rect 25468 -11300 27930 -11248
rect 25468 -12096 25552 -11300
rect 26182 -12096 27930 -11300
rect 25468 -12176 27930 -12096
rect -582 -16188 40 -16174
rect -13502 -16808 40 -16188
rect -13502 -17200 -1018 -16808
rect -574 -17200 40 -16808
rect -13502 -17242 40 -17200
rect -13502 -17304 38 -17242
rect -13502 -17400 -202 -17304
rect -6682 -18522 -5352 -18382
rect -6682 -19054 -6384 -18522
rect -5662 -19054 -5352 -18522
rect -22160 -20188 -21434 -19764
rect -22164 -20682 -21224 -20188
rect -6682 -20342 -5352 -19054
use dac_cell1  dac_cell1_0
timestamp 1697955996
transform 1 0 -1148 0 1 8720
box -3902 -1834 10992 3012
use dac_cell2  dac_cell2_0
timestamp 1697955996
transform 1 0 -2028 0 1 -378
box -3290 40 5010 5340
use dac_cell3  dac_cell3_0
timestamp 1697955996
transform 1 0 1882 0 1 -5798
box -4704 -2118 1052 4150
use dac_cell4  dac_cell4_0
timestamp 1697955996
transform 1 0 -1562 0 1 -15346
box -278 -1932 4578 5878
use esd_structure  esd_structure_0
timestamp 1698216219
transform 1 0 -16808 0 1 -2800
box -4892 -2846 654 2614
use esd_structure  esd_structure_1
timestamp 1698216219
transform 1 0 -16856 0 1 8610
box -4892 -2846 654 2614
use esd_structure  esd_structure_2
timestamp 1698216219
transform 1 0 -16808 0 1 2850
box -4892 -2846 654 2614
use esd_structure  esd_structure_3
timestamp 1698216219
transform -1 0 16354 0 -1 -11734
box -4892 -2846 654 2614
use esd_structure  esd_structure_4
timestamp 1698216219
transform 1 0 -16808 0 1 -8490
box -4892 -2846 654 2614
use esd_structure  esd_structure_5
timestamp 1698216219
transform 1 0 -16758 0 1 -14100
box -4892 -2846 654 2614
use miel21_opamp  miel21_opamp_0
timestamp 1697955996
transform 1 0 12484 0 1 -6200
box -3496 2114 9690 10290
use sky130_fd_pr__res_high_po_5p73_6QQPRG  sky130_fd_pr__res_high_po_5p73_6QQPRG_0
timestamp 1697955996
transform 0 1 -9495 -1 0 -13405
box -739 -723 739 723
use sky130_fd_pr__res_high_po_5p73_6QQPRG  sky130_fd_pr__res_high_po_5p73_6QQPRG_1
timestamp 1697955996
transform 0 1 -9505 -1 0 -14867
box -739 -723 739 723
use sky130_fd_pr__res_high_po_5p73_6QQPRG  sky130_fd_pr__res_high_po_5p73_6QQPRG_2
timestamp 1697955996
transform 0 1 -9517 -1 0 -16361
box -739 -723 739 723
use sky130_fd_pr__res_xhigh_po_0p35_PZAK34  sky130_fd_pr__res_xhigh_po_0p35_PZAK34_0
timestamp 1697955996
transform 0 1 16306 -1 0 6255
box -201 -1018 201 1018
use sky130_fd_pr__res_xhigh_po_0p35_PZAK34  sky130_fd_pr__res_xhigh_po_0p35_PZAK34_1
timestamp 1697955996
transform 0 1 16316 -1 0 5815
box -201 -1018 201 1018
use sky130_fd_pr__res_xhigh_po_0p35_PZAK34  sky130_fd_pr__res_xhigh_po_0p35_PZAK34_2
timestamp 1697955996
transform 0 1 16296 -1 0 6683
box -201 -1018 201 1018
use sky130_fd_pr__res_xhigh_po_2p85_5DPYAB  sky130_fd_pr__res_xhigh_po_2p85_5DPYAB_0
timestamp 1697955996
transform 0 1 8741 -1 0 -10857
box -451 -723 451 723
use sky130_fd_pr__res_xhigh_po_2p85_5DPYAB  sky130_fd_pr__res_xhigh_po_2p85_5DPYAB_1
timestamp 1697955996
transform 0 1 8753 -1 0 -9063
box -451 -723 451 723
use sky130_fd_pr__res_xhigh_po_2p85_5DPYAB  sky130_fd_pr__res_xhigh_po_2p85_5DPYAB_2
timestamp 1697955996
transform 0 1 8737 -1 0 -11757
box -451 -723 451 723
use sky130_fd_pr__res_high_po_5p73_6QQPRG  XR1
timestamp 1697955996
transform 0 1 -9539 -1 0 -17825
box -739 -723 739 723
use sky130_fd_pr__res_xhigh_po_2p85_5DPYAB  XR2
timestamp 1697955996
transform 0 1 8747 -1 0 -9957
box -451 -723 451 723
use sky130_fd_pr__res_xhigh_po_0p35_PZAK34  XR3
timestamp 1697955996
transform 0 1 16304 -1 0 5395
box -201 -1018 201 1018
<< labels >>
rlabel metal1 7054 -334 7314 894 1 op_amp_in
rlabel metal1 -8412 -14134 -8106 -13372 1 in_iref
flabel metal3 -6420 -20098 -6220 -19898 0 FreeSans 1280 0 0 0 vgnd
port 5 nsew
flabel metal3 -4850 13056 -4650 13256 0 FreeSans 1280 0 0 0 vsup
port 6 nsew
flabel metal3 25188 -168 25388 32 0 FreeSans 1280 0 0 0 out
port 7 nsew
flabel metal3 26818 -11864 27018 -11664 0 FreeSans 1280 0 0 0 vbias18
port 8 nsew
flabel metal3 -27704 8550 -27504 8750 0 FreeSans 1280 0 0 0 in1
port 0 nsew
flabel metal3 -27480 2688 -27280 2888 0 FreeSans 1280 0 0 0 in2
port 1 nsew
flabel metal3 -27482 -3166 -27282 -2966 0 FreeSans 1280 0 0 0 in3
port 2 nsew
flabel metal3 -27444 -8652 -27244 -8452 0 FreeSans 1280 0 0 0 in4
port 3 nsew
flabel metal3 -21726 -20602 -21526 -20402 0 FreeSans 1280 0 0 0 vbias07
port 4 nsew
rlabel metal2 -6520 -15434 -6174 -13688 1 vbias_v
<< end >>
