magic
tech sky130A
timestamp 1697384985
<< nwell >>
rect -179 -198 179 198
<< mvpmos >>
rect -50 -50 50 50
<< mvpdiff >>
rect -79 44 -50 50
rect -79 -44 -73 44
rect -56 -44 -50 44
rect -79 -50 -50 -44
rect 50 44 79 50
rect 50 -44 56 44
rect 73 -44 79 44
rect 50 -50 79 -44
<< mvpdiffc >>
rect -73 -44 -56 44
rect 56 -44 73 44
<< mvnsubdiff >>
rect -146 159 146 165
rect -146 142 -92 159
rect 92 142 146 159
rect -146 136 146 142
rect -146 111 -117 136
rect -146 -111 -140 111
rect -123 -111 -117 111
rect 117 111 146 136
rect -146 -136 -117 -111
rect 117 -111 123 111
rect 140 -111 146 111
rect 117 -136 146 -111
rect -146 -142 146 -136
rect -146 -159 -92 -142
rect 92 -159 146 -142
rect -146 -165 146 -159
<< mvnsubdiffcont >>
rect -92 142 92 159
rect -140 -111 -123 111
rect 123 -111 140 111
rect -92 -159 92 -142
<< poly >>
rect -50 90 50 98
rect -50 73 -42 90
rect 42 73 50 90
rect -50 50 50 73
rect -50 -73 50 -50
rect -50 -90 -42 -73
rect 42 -90 50 -73
rect -50 -98 50 -90
<< polycont >>
rect -42 73 42 90
rect -42 -90 42 -73
<< locali >>
rect -140 142 -92 159
rect 92 142 140 159
rect -140 111 -123 142
rect 123 111 140 142
rect -50 73 -42 90
rect 42 73 50 90
rect -73 44 -56 52
rect -73 -52 -56 -44
rect 56 44 73 52
rect 56 -52 73 -44
rect -50 -90 -42 -73
rect 42 -90 50 -73
rect -140 -142 -123 -111
rect 123 -142 140 -111
rect -140 -159 -92 -142
rect 92 -159 140 -142
<< viali >>
rect -42 73 42 90
rect -73 -44 -56 44
rect 56 -44 73 44
rect -42 -90 42 -73
<< metal1 >>
rect -48 90 48 93
rect -48 73 -42 90
rect 42 73 48 90
rect -48 70 48 73
rect -76 44 -53 50
rect -76 -44 -73 44
rect -56 -44 -53 44
rect -76 -50 -53 -44
rect 53 44 76 50
rect 53 -44 56 44
rect 73 -44 76 44
rect 53 -50 76 -44
rect -48 -73 48 -70
rect -48 -90 -42 -73
rect 42 -90 48 -73
rect -48 -93 48 -90
<< properties >>
string FIXED_BBOX -131 -151 131 151
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
