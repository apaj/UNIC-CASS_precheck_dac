**.subckt dIV05
D1 out GND sky130_fd_pr__diode_pw2nd_05v5 area=1e+12
V1 in GND 3
R1 out in 1k m=1
**** begin user architecture code


.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.param mc_pr_switch=0
*** ANALYSIS TO DO
.dc V1 -5 5 0.01

.control
set wr_vecnames
set wr_singlescale
run
******** results filename  ************ nodes to write
save in out i(V1)
plot 0-i(V1)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
