magic
tech sky130A
magscale 1 2
timestamp 1697704145
<< nwell >>
rect -358 -1097 358 1097
<< mvpmos >>
rect -100 -800 100 800
<< mvpdiff >>
rect -158 788 -100 800
rect -158 -788 -146 788
rect -112 -788 -100 788
rect -158 -800 -100 -788
rect 100 788 158 800
rect 100 -788 112 788
rect 146 -788 158 788
rect 100 -800 158 -788
<< mvpdiffc >>
rect -146 -788 -112 788
rect 112 -788 146 788
<< mvnsubdiff >>
rect -292 1019 292 1031
rect -292 985 -184 1019
rect 184 985 292 1019
rect -292 973 292 985
rect -292 923 -234 973
rect -292 -923 -280 923
rect -246 -923 -234 923
rect 234 923 292 973
rect -292 -973 -234 -923
rect 234 -923 246 923
rect 280 -923 292 923
rect 234 -973 292 -923
rect -292 -985 292 -973
rect -292 -1019 -184 -985
rect 184 -1019 292 -985
rect -292 -1031 292 -1019
<< mvnsubdiffcont >>
rect -184 985 184 1019
rect -280 -923 -246 923
rect 246 -923 280 923
rect -184 -1019 184 -985
<< poly >>
rect -100 881 100 897
rect -100 847 -84 881
rect 84 847 100 881
rect -100 800 100 847
rect -100 -847 100 -800
rect -100 -881 -84 -847
rect 84 -881 100 -847
rect -100 -897 100 -881
<< polycont >>
rect -84 847 84 881
rect -84 -881 84 -847
<< locali >>
rect -280 985 -184 1019
rect 184 985 280 1019
rect -280 923 -246 985
rect 246 923 280 985
rect -100 847 -84 881
rect 84 847 100 881
rect -146 788 -112 804
rect -146 -804 -112 -788
rect 112 788 146 804
rect 112 -804 146 -788
rect -100 -881 -84 -847
rect 84 -881 100 -847
rect -280 -985 -246 -923
rect 246 -985 280 -923
rect -280 -1019 -184 -985
rect 184 -1019 280 -985
<< viali >>
rect -84 847 84 881
rect -146 -788 -112 788
rect 112 -788 146 788
rect -84 -881 84 -847
<< metal1 >>
rect -96 881 96 887
rect -96 847 -84 881
rect 84 847 96 881
rect -96 841 96 847
rect -152 788 -106 800
rect -152 -788 -146 788
rect -112 -788 -106 788
rect -152 -800 -106 -788
rect 106 788 152 800
rect 106 -788 112 788
rect 146 -788 152 788
rect 106 -800 152 -788
rect -96 -847 96 -841
rect -96 -881 -84 -847
rect 84 -881 96 -847
rect -96 -887 96 -881
<< properties >>
string FIXED_BBOX -263 -1002 263 1002
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 8.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
