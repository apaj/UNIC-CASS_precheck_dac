* SPICE3 file created from dac_cell1.ext - technology: sky130A

.option scale=5000u

.subckt dac_cell1 vsup vgnd iref vsw iout iout_n vbias
X0 m1_10330_1196# vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=11600
X1 m1_10330_1196# vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=11600
X2 m1_10330_1196# vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=11600
X3 m1_10330_1196# vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=11600
X4 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 ad=11600 pd=516 as=23200 ps=1032 w=200 l=200
X5 li_n800_n926# iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X6 iout vsw li_n800_n926# vsup sky130_fd_pr__pfet_g5v0d10v5 ad=11600 pd=516 as=0 ps=0 w=200 l=200
X7 iout_n vbias li_n800_n926# vsup sky130_fd_pr__pfet_g5v0d10v5 ad=11600 pd=516 as=0 ps=0 w=200 l=200
.ends
