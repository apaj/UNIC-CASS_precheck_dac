magic
tech sky130A
timestamp 1698258108
use dac_top_cell  dac_top_cell_0
timestamp 1698257525
transform 1 0 12271 0 1 9577
box -14014 -10341 13965 9172
<< end >>
