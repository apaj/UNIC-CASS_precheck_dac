**.subckt tb_dac_top_cell_tran
vsw1 vsw1 GND pulse(0, 3.3, 20ms, 1ns, 1ns, 10ms, 20ms)
vsw2 vsw2 GND pulse(0, 3.3, 20ms, 1ns, 1ns, 20ms, 40ms)
vsw3 vsw3 GND pulse(0, 3.3, 20ms, 1ns, 1ns, 40ms, 80ms)
vsw4 vsw4 GND pulse(0, 3.3, 20ms, 1ns, 1ns, 80ms, 160ms)
Rout1 vout GND 1k m=1
Vsup net1 GND 3.3
Vbias07 net2 GND 0.7
x1 vsw1 vsw2 vsw3 vout vsw4 net3 net2 net1 GND dac_top_cell
Vbias18 net3 GND 1.8
**** begin user architecture code


.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.param mc_pr_switch=0
*** ANALYSIS TO DO

.tran 0.1 500m 0.001m
.save vout
.save x1.op_amp_in
.save vsw1 vsw2 vsw3 vsw4

.control
set wr_vecnames
set wr_singlescale

run
******** results filename  ************ nodes to write
wrdata $DEV_PATH/res/dac_top_cell_vout_tran_vol.res vout
wrdata $DEV_PATH/res/dac_top_cell_vsw1_tran_vol.res vsw1
wrdata $DEV_PATH/res/dac_top_cell_vsw2_tran_vol.res vsw2
wrdata $DEV_PATH/res/dac_top_cell_vsw3_tran_vol.res vsw3
wrdata $DEV_PATH/res/dac_top_cell_vsw4_tran_vol.res vsw4
.endc


**** end user architecture code
**.ends

* expanding   symbol:  dac_top_cell.sym # of pins=9
* sym_path: /opt/uniccass/dev/top_cell_esd/tb/dac_top_cell.sym
* sch_path: /opt/uniccass/dev/top_cell_esd/tb/dac_top_cell.sch
.subckt dac_top_cell  in1 in2 in3 out in4 vbias18 vbias07 vsup vgnd
*.iopin in1
*.iopin in2
*.iopin in3
*.iopin in4
*.iopin vbias07
*.iopin vgnd
*.iopin vsup
*.iopin out
*.iopin vbias18
x2 vsup in_iref vgnd net2 vbias_v net5 vgnd dac_cell2
x3 vsup vgnd in_iref net3 vbias_v net5 vgnd dac_cell3
x4 vsup in_iref vgnd net4 vbias_v net5 vgnd dac_cell4
x5 vsup out op_amp_in net9 vgnd miel21_opamp
x1 vsup in_iref vgnd net1 vbias_v net5 vgnd dac_cell1
XR1 net6 net5 vgnd sky130_fd_pr__res_xhigh_po_2p85 L=1.25 mult=1 m=1
XR2 op_amp_in net6 vgnd sky130_fd_pr__res_xhigh_po_2p85 L=1.25 mult=1 m=1
XR4 net6 net5 vgnd sky130_fd_pr__res_xhigh_po_2p85 L=1.25 mult=1 m=1
XR3 op_amp_in net6 vgnd sky130_fd_pr__res_xhigh_po_2p85 L=1.25 mult=1 m=1
XR5 net7 op_amp_in vgnd sky130_fd_pr__res_xhigh_po_0p35 L=4.2 mult=1 m=1
XR6 out net7 vgnd sky130_fd_pr__res_xhigh_po_0p35 L=4.2 mult=1 m=1
XR7 net7 op_amp_in vgnd sky130_fd_pr__res_xhigh_po_0p35 L=4.2 mult=1 m=1
XR8 out net7 vgnd sky130_fd_pr__res_xhigh_po_0p35 L=4.2 mult=1 m=1
XR9 net8 in_iref vgnd sky130_fd_pr__res_high_po_5p73 L=1.25 mult=1 m=1
XR10 net8 in_iref vgnd sky130_fd_pr__res_high_po_5p73 L=1.25 mult=1 m=1
XR11 vgnd net8 vgnd sky130_fd_pr__res_high_po_5p73 L=1.25 mult=1 m=1
XR12 vgnd net8 vgnd sky130_fd_pr__res_high_po_5p73 L=1.25 mult=1 m=1
x6 vsup in1 net1 vgnd esd_cell
x7 vsup in2 net2 vgnd esd_cell
x8 vsup in3 net3 vgnd esd_cell
x9 vsup in4 net4 vgnd esd_cell
x10 vsup vbias07 vbias_v vgnd esd_cell
x11 vsup vbias18 net9 vgnd esd_cell
.ends


* expanding   symbol:  /opt/uniccass/dev/dac_cell2/tb/dac_cell2.sym # of pins=7
* sym_path: /opt/uniccass/dev/dac_cell2/tb/dac_cell2.sym
* sch_path: /opt/uniccass/dev/dac_cell2/tb/dac_cell2.sch
.subckt dac_cell2  vsup iref vgnd vsw vbias iout_n iout
*.iopin vsup
*.iopin vgnd
*.iopin iref
*.iopin vsw
*.iopin iout
*.iopin iout_n
*.iopin vbias
XM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 sourceM3M4 iref sourceM2 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 iout vsw sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 iout_n vbias sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XR1 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=1 m=1
XR2 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=1 m=1
XR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=1 m=1
XR4 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=1 m=1
.ends


* expanding   symbol:  /opt/uniccass/dev/dac_cell3/tb/dac_cell3.sym # of pins=7
* sym_path: /opt/uniccass/dev/dac_cell3/tb/dac_cell3.sym
* sch_path: /opt/uniccass/dev/dac_cell3/tb/dac_cell3.sch
.subckt dac_cell3  vsup vgnd iref vsw vbias iout_n iout
*.iopin vsup
*.iopin vgnd
*.iopin iref
*.iopin vsw
*.iopin iout
*.iopin iout_n
*.iopin vbias
XM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 sourceM3M4 iref sourceM2 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 iout vsw sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 iout_n vbias sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XR1 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR2 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR4 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
.ends


* expanding   symbol:  /opt/uniccass/dev/dac_cell4/tb/dac_cell4.sym # of pins=7
* sym_path: /opt/uniccass/dev/dac_cell4/tb/dac_cell4.sym
* sch_path: /opt/uniccass/dev/dac_cell4/tb/dac_cell4.sch
.subckt dac_cell4  vsup iref vgnd vsw vbias iout_n iout
*.iopin vsup
*.iopin vgnd
*.iopin iref
*.iopin vsw
*.iopin iout
*.iopin iout_n
*.iopin vbias
XM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 sourceM3M4 iref sourceM2 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 iout vsw sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 iout_n vbias sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XR1 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=6.3 mult=1 m=1
XR2 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=6.3 mult=1 m=1
XR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=6.3 mult=1 m=1
XR4 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=6.3 mult=1 m=1
.ends


* expanding   symbol:  /opt/uniccass/dev/opamp/miel21_opamp.sym # of pins=5
* sym_path: /opt/uniccass/dev/opamp/miel21_opamp.sym
* sch_path: /opt/uniccass/dev/opamp/miel21_opamp.sch
.subckt miel21_opamp  power outSingle inPos inNeg ground
*.ipin inPos
*.ipin inNeg
*.opin outSingle
*.iopin power
*.iopin ground
XM6 d1 d1 power power sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=21 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 d2 d1 power power sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=21 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 outSingle d2 power power sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=100 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM1 d1 inPos nsources ground sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM2 d2 inNeg nsources ground sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 bias bias ground ground sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 nsources bias ground ground sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM5 outSingle bias ground ground sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=48 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XR1 bias net2 ground sky130_fd_pr__res_xhigh_po_0p69 L=6 mult=1 m=1
XC1 outSingle d2 sky130_fd_pr__cap_mim_m3_1 W=10 L=14 MF=1 m=1
XR2 net2 net1 ground sky130_fd_pr__res_xhigh_po_0p69 L=6 mult=1 m=1
XR3 net1 power ground sky130_fd_pr__res_xhigh_po_0p69 L=6 mult=1 m=1
.ends


* expanding   symbol:  /opt/uniccass/dev/dac_cell1/tb/dac_cell1.sym # of pins=7
* sym_path: /opt/uniccass/dev/dac_cell1/tb/dac_cell1.sym
* sch_path: /opt/uniccass/dev/dac_cell1/tb/dac_cell1.sch
.subckt dac_cell1  vsup iref vgnd vsw vbias iout_n iout
*.iopin vsup
*.iopin vgnd
*.iopin iref
*.iopin vsw
*.iopin iout
*.iopin iout_n
*.iopin vbias
XM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 sourceM3M4 iref sourceM2 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 iout vsw sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 iout_n vbias sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XR1 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
XR2 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
XR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
XR4 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
.ends


* expanding   symbol:  /opt/uniccass/dev/esd_cell/tb/esd_cell.sym # of pins=4
* sym_path: /opt/uniccass/dev/esd_cell/tb/esd_cell.sym
* sch_path: /opt/uniccass/dev/esd_cell/tb/esd_cell.sch
.subckt esd_cell  vsup pad gate vgnd
*.iopin vsup
*.iopin pad
*.iopin vgnd
*.iopin gate
D1 pad vsup sky130_fd_pr__diode_pd2nw_11v0 area=10e+18
D3 gate vsup sky130_fd_pr__diode_pd2nw_05v5 area=0.203e+18
D4 vgnd gate sky130_fd_pr__diode_pw2nd_05v5 area=0.203e+18
XR1 gate pad vgnd sky130_fd_pr__res_high_po W=0.35 L=10 mult=1 m=1
D8 vgnd pad sky130_fd_pr__diode_pw2nd_11v0 area=10e+18
D2 pad vsup sky130_fd_pr__diode_pd2nw_11v0 area=10e+18
D5 pad vsup sky130_fd_pr__diode_pd2nw_11v0 area=10e+18
D6 pad vsup sky130_fd_pr__diode_pd2nw_11v0 area=10e+18
D7 pad vsup sky130_fd_pr__diode_pd2nw_11v0 area=10e+18
D9 vgnd pad sky130_fd_pr__diode_pw2nd_11v0 area=10e+18
D10 vgnd pad sky130_fd_pr__diode_pw2nd_11v0 area=10e+18
D11 vgnd pad sky130_fd_pr__diode_pw2nd_11v0 area=10e+18
D12 vgnd pad sky130_fd_pr__diode_pw2nd_11v0 area=10e+18
.ends

.GLOBAL GND
** flattened .save nodes
.save vout
.save x1.op_amp_in
.save vsw1 vsw2 vsw3 vsw4
.end
