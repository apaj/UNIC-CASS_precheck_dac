magic
tech sky130A
magscale 1 2
timestamp 1695142129
<< dnwell >>
rect -876 -5937 876 5937
<< nwell >>
rect -956 5731 956 6017
rect -956 -5731 -670 5731
rect 670 -5731 956 5731
rect -956 -6017 956 -5731
<< pwell >>
rect -670 5573 -140 5731
rect -670 115 -140 273
rect 140 5573 670 5731
rect 140 115 670 273
rect -670 -273 -140 -115
rect -670 -5731 -140 -5573
rect 140 -273 670 -115
rect 140 -5731 670 -5573
<< rpw >>
rect -670 273 -140 5573
rect 140 273 670 5573
rect -670 -5573 -140 -273
rect 140 -5573 670 -273
<< psubdiff >>
rect -630 5573 -606 5679
rect -204 5573 -180 5679
rect 180 5573 204 5679
rect 606 5573 630 5679
rect -630 167 -606 273
rect -204 167 -180 273
rect 180 167 204 273
rect 606 167 630 273
rect -630 -273 -606 -167
rect -204 -273 -180 -167
rect 180 -273 204 -167
rect 606 -273 630 -167
rect -630 -5679 -606 -5573
rect -204 -5679 -180 -5573
rect 180 -5679 204 -5573
rect 606 -5679 630 -5573
<< nsubdiff >>
rect -830 5857 -734 5891
rect 734 5857 830 5891
rect -830 5795 -796 5857
rect 796 5795 830 5857
rect -830 -5857 -796 -5795
rect 796 -5857 830 -5795
rect -830 -5891 -734 -5857
rect 734 -5891 830 -5857
<< psubdiffcont >>
rect -606 5573 -204 5679
rect 204 5573 606 5679
rect -606 167 -204 273
rect 204 167 606 273
rect -606 -273 -204 -167
rect 204 -273 606 -167
rect -606 -5679 -204 -5573
rect 204 -5679 606 -5573
<< nsubdiffcont >>
rect -734 5857 734 5891
rect -830 -5795 -796 5795
rect 796 -5795 830 5795
rect -734 -5891 734 -5857
<< locali >>
rect -830 5857 -734 5891
rect 734 5857 830 5891
rect -830 5795 -796 5857
rect 796 5795 830 5857
rect -622 5643 -606 5679
rect -204 5643 -188 5679
rect -622 5590 -618 5643
rect -192 5590 -188 5643
rect -622 5573 -606 5590
rect -204 5573 -188 5590
rect 188 5643 204 5679
rect 606 5643 622 5679
rect 188 5590 192 5643
rect 618 5590 622 5643
rect 188 5573 204 5590
rect 606 5573 622 5590
rect -622 256 -606 273
rect -204 256 -188 273
rect -622 203 -618 256
rect -192 203 -188 256
rect -622 167 -606 203
rect -204 167 -188 203
rect 188 256 204 273
rect 606 256 622 273
rect 188 203 192 256
rect 618 203 622 256
rect 188 167 204 203
rect 606 167 622 203
rect -622 -203 -606 -167
rect -204 -203 -188 -167
rect -622 -256 -618 -203
rect -192 -256 -188 -203
rect -622 -273 -606 -256
rect -204 -273 -188 -256
rect 188 -203 204 -167
rect 606 -203 622 -167
rect 188 -256 192 -203
rect 618 -256 622 -203
rect 188 -273 204 -256
rect 606 -273 622 -256
rect -622 -5590 -606 -5573
rect -204 -5590 -188 -5573
rect -622 -5643 -618 -5590
rect -192 -5643 -188 -5590
rect -622 -5679 -606 -5643
rect -204 -5679 -188 -5643
rect 188 -5590 204 -5573
rect 606 -5590 622 -5573
rect 188 -5643 192 -5590
rect 618 -5643 622 -5590
rect 188 -5679 204 -5643
rect 606 -5679 622 -5643
rect -830 -5857 -796 -5795
rect 796 -5857 830 -5795
rect -830 -5891 -734 -5857
rect 734 -5891 830 -5857
<< viali >>
rect -618 5590 -606 5643
rect -606 5590 -204 5643
rect -204 5590 -192 5643
rect 192 5590 204 5643
rect 204 5590 606 5643
rect 606 5590 618 5643
rect -618 203 -606 256
rect -606 203 -204 256
rect -204 203 -192 256
rect 192 203 204 256
rect 204 203 606 256
rect 606 203 618 256
rect -618 -256 -606 -203
rect -606 -256 -204 -203
rect -204 -256 -192 -203
rect 192 -256 204 -203
rect 204 -256 606 -203
rect 606 -256 618 -203
rect -618 -5643 -606 -5590
rect -606 -5643 -204 -5590
rect -204 -5643 -192 -5590
rect 192 -5643 204 -5590
rect 204 -5643 606 -5590
rect 606 -5643 618 -5590
<< metal1 >>
rect -630 5643 -180 5649
rect -630 5590 -618 5643
rect -192 5590 -180 5643
rect -630 5584 -180 5590
rect 180 5643 630 5649
rect 180 5590 192 5643
rect 618 5590 630 5643
rect 180 5584 630 5590
rect -630 256 -180 262
rect -630 203 -618 256
rect -192 203 -180 256
rect -630 197 -180 203
rect 180 256 630 262
rect 180 203 192 256
rect 618 203 630 256
rect 180 197 630 203
rect -630 -203 -180 -197
rect -630 -256 -618 -203
rect -192 -256 -180 -203
rect -630 -262 -180 -256
rect 180 -203 630 -197
rect 180 -256 192 -203
rect 618 -256 630 -203
rect 180 -262 630 -256
rect -630 -5590 -180 -5584
rect -630 -5643 -618 -5590
rect -192 -5643 -180 -5590
rect -630 -5649 -180 -5643
rect 180 -5590 630 -5584
rect 180 -5643 192 -5590
rect 618 -5643 630 -5590
rect 180 -5649 630 -5643
<< properties >>
string FIXED_BBOX -813 -5874 813 5874
string gencell sky130_fd_pr__res_iso_pw
string library sky130
string parameters w 2.650 l 26.50 m 2 nx 2 wmin 2.650 lmin 26.50 rho 975 val 10.766k dummy 0 dw 0.25 term 1.0 guard 1 endcov 100 full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
