magic
tech sky130A
magscale 1 2
timestamp 1697933062
<< pwell >>
rect -1251 -858 1251 858
<< mvnmos >>
rect -1023 -600 -923 600
rect -745 -600 -645 600
rect -467 -600 -367 600
rect -189 -600 -89 600
rect 89 -600 189 600
rect 367 -600 467 600
rect 645 -600 745 600
rect 923 -600 1023 600
<< mvndiff >>
rect -1081 588 -1023 600
rect -1081 -588 -1069 588
rect -1035 -588 -1023 588
rect -1081 -600 -1023 -588
rect -923 588 -865 600
rect -923 -588 -911 588
rect -877 -588 -865 588
rect -923 -600 -865 -588
rect -803 588 -745 600
rect -803 -588 -791 588
rect -757 -588 -745 588
rect -803 -600 -745 -588
rect -645 588 -587 600
rect -645 -588 -633 588
rect -599 -588 -587 588
rect -645 -600 -587 -588
rect -525 588 -467 600
rect -525 -588 -513 588
rect -479 -588 -467 588
rect -525 -600 -467 -588
rect -367 588 -309 600
rect -367 -588 -355 588
rect -321 -588 -309 588
rect -367 -600 -309 -588
rect -247 588 -189 600
rect -247 -588 -235 588
rect -201 -588 -189 588
rect -247 -600 -189 -588
rect -89 588 -31 600
rect -89 -588 -77 588
rect -43 -588 -31 588
rect -89 -600 -31 -588
rect 31 588 89 600
rect 31 -588 43 588
rect 77 -588 89 588
rect 31 -600 89 -588
rect 189 588 247 600
rect 189 -588 201 588
rect 235 -588 247 588
rect 189 -600 247 -588
rect 309 588 367 600
rect 309 -588 321 588
rect 355 -588 367 588
rect 309 -600 367 -588
rect 467 588 525 600
rect 467 -588 479 588
rect 513 -588 525 588
rect 467 -600 525 -588
rect 587 588 645 600
rect 587 -588 599 588
rect 633 -588 645 588
rect 587 -600 645 -588
rect 745 588 803 600
rect 745 -588 757 588
rect 791 -588 803 588
rect 745 -600 803 -588
rect 865 588 923 600
rect 865 -588 877 588
rect 911 -588 923 588
rect 865 -600 923 -588
rect 1023 588 1081 600
rect 1023 -588 1035 588
rect 1069 -588 1081 588
rect 1023 -600 1081 -588
<< mvndiffc >>
rect -1069 -588 -1035 588
rect -911 -588 -877 588
rect -791 -588 -757 588
rect -633 -588 -599 588
rect -513 -588 -479 588
rect -355 -588 -321 588
rect -235 -588 -201 588
rect -77 -588 -43 588
rect 43 -588 77 588
rect 201 -588 235 588
rect 321 -588 355 588
rect 479 -588 513 588
rect 599 -588 633 588
rect 757 -588 791 588
rect 877 -588 911 588
rect 1035 -588 1069 588
<< mvpsubdiff >>
rect -1215 810 1215 822
rect -1215 776 -1107 810
rect 1107 776 1215 810
rect -1215 764 1215 776
rect -1215 714 -1157 764
rect -1215 -714 -1203 714
rect -1169 -714 -1157 714
rect 1157 714 1215 764
rect -1215 -764 -1157 -714
rect 1157 -714 1169 714
rect 1203 -714 1215 714
rect 1157 -764 1215 -714
rect -1215 -776 1215 -764
rect -1215 -810 -1107 -776
rect 1107 -810 1215 -776
rect -1215 -822 1215 -810
<< mvpsubdiffcont >>
rect -1107 776 1107 810
rect -1203 -714 -1169 714
rect 1169 -714 1203 714
rect -1107 -810 1107 -776
<< poly >>
rect -1023 672 -923 688
rect -1023 638 -1007 672
rect -939 638 -923 672
rect -1023 600 -923 638
rect -745 672 -645 688
rect -745 638 -729 672
rect -661 638 -645 672
rect -745 600 -645 638
rect -467 672 -367 688
rect -467 638 -451 672
rect -383 638 -367 672
rect -467 600 -367 638
rect -189 672 -89 688
rect -189 638 -173 672
rect -105 638 -89 672
rect -189 600 -89 638
rect 89 672 189 688
rect 89 638 105 672
rect 173 638 189 672
rect 89 600 189 638
rect 367 672 467 688
rect 367 638 383 672
rect 451 638 467 672
rect 367 600 467 638
rect 645 672 745 688
rect 645 638 661 672
rect 729 638 745 672
rect 645 600 745 638
rect 923 672 1023 688
rect 923 638 939 672
rect 1007 638 1023 672
rect 923 600 1023 638
rect -1023 -638 -923 -600
rect -1023 -672 -1007 -638
rect -939 -672 -923 -638
rect -1023 -688 -923 -672
rect -745 -638 -645 -600
rect -745 -672 -729 -638
rect -661 -672 -645 -638
rect -745 -688 -645 -672
rect -467 -638 -367 -600
rect -467 -672 -451 -638
rect -383 -672 -367 -638
rect -467 -688 -367 -672
rect -189 -638 -89 -600
rect -189 -672 -173 -638
rect -105 -672 -89 -638
rect -189 -688 -89 -672
rect 89 -638 189 -600
rect 89 -672 105 -638
rect 173 -672 189 -638
rect 89 -688 189 -672
rect 367 -638 467 -600
rect 367 -672 383 -638
rect 451 -672 467 -638
rect 367 -688 467 -672
rect 645 -638 745 -600
rect 645 -672 661 -638
rect 729 -672 745 -638
rect 645 -688 745 -672
rect 923 -638 1023 -600
rect 923 -672 939 -638
rect 1007 -672 1023 -638
rect 923 -688 1023 -672
<< polycont >>
rect -1007 638 -939 672
rect -729 638 -661 672
rect -451 638 -383 672
rect -173 638 -105 672
rect 105 638 173 672
rect 383 638 451 672
rect 661 638 729 672
rect 939 638 1007 672
rect -1007 -672 -939 -638
rect -729 -672 -661 -638
rect -451 -672 -383 -638
rect -173 -672 -105 -638
rect 105 -672 173 -638
rect 383 -672 451 -638
rect 661 -672 729 -638
rect 939 -672 1007 -638
<< locali >>
rect -1203 776 -1107 810
rect 1107 776 1203 810
rect -1203 714 -1169 776
rect 1169 714 1203 776
rect -1023 638 -1007 672
rect -939 638 -923 672
rect -745 638 -729 672
rect -661 638 -645 672
rect -467 638 -451 672
rect -383 638 -367 672
rect -189 638 -173 672
rect -105 638 -89 672
rect 89 638 105 672
rect 173 638 189 672
rect 367 638 383 672
rect 451 638 467 672
rect 645 638 661 672
rect 729 638 745 672
rect 923 638 939 672
rect 1007 638 1023 672
rect -1069 588 -1035 604
rect -1069 -604 -1035 -588
rect -911 588 -877 604
rect -911 -604 -877 -588
rect -791 588 -757 604
rect -791 -604 -757 -588
rect -633 588 -599 604
rect -633 -604 -599 -588
rect -513 588 -479 604
rect -513 -604 -479 -588
rect -355 588 -321 604
rect -355 -604 -321 -588
rect -235 588 -201 604
rect -235 -604 -201 -588
rect -77 588 -43 604
rect -77 -604 -43 -588
rect 43 588 77 604
rect 43 -604 77 -588
rect 201 588 235 604
rect 201 -604 235 -588
rect 321 588 355 604
rect 321 -604 355 -588
rect 479 588 513 604
rect 479 -604 513 -588
rect 599 588 633 604
rect 599 -604 633 -588
rect 757 588 791 604
rect 757 -604 791 -588
rect 877 588 911 604
rect 877 -604 911 -588
rect 1035 588 1069 604
rect 1035 -604 1069 -588
rect -1023 -672 -1007 -638
rect -939 -672 -923 -638
rect -745 -672 -729 -638
rect -661 -672 -645 -638
rect -467 -672 -451 -638
rect -383 -672 -367 -638
rect -189 -672 -173 -638
rect -105 -672 -89 -638
rect 89 -672 105 -638
rect 173 -672 189 -638
rect 367 -672 383 -638
rect 451 -672 467 -638
rect 645 -672 661 -638
rect 729 -672 745 -638
rect 923 -672 939 -638
rect 1007 -672 1023 -638
rect -1203 -776 -1169 -714
rect 1169 -776 1203 -714
rect -1203 -810 -1107 -776
rect 1107 -810 1203 -776
<< viali >>
rect -1007 638 -939 672
rect -729 638 -661 672
rect -451 638 -383 672
rect -173 638 -105 672
rect 105 638 173 672
rect 383 638 451 672
rect 661 638 729 672
rect 939 638 1007 672
rect -1069 -588 -1035 588
rect -911 -588 -877 588
rect -791 -588 -757 588
rect -633 -588 -599 588
rect -513 -588 -479 588
rect -355 -588 -321 588
rect -235 -588 -201 588
rect -77 -588 -43 588
rect 43 -588 77 588
rect 201 -588 235 588
rect 321 -588 355 588
rect 479 -588 513 588
rect 599 -588 633 588
rect 757 -588 791 588
rect 877 -588 911 588
rect 1035 -588 1069 588
rect -1007 -672 -939 -638
rect -729 -672 -661 -638
rect -451 -672 -383 -638
rect -173 -672 -105 -638
rect 105 -672 173 -638
rect 383 -672 451 -638
rect 661 -672 729 -638
rect 939 -672 1007 -638
<< metal1 >>
rect -1019 672 -927 678
rect -1019 638 -1007 672
rect -939 638 -927 672
rect -1019 632 -927 638
rect -741 672 -649 678
rect -741 638 -729 672
rect -661 638 -649 672
rect -741 632 -649 638
rect -463 672 -371 678
rect -463 638 -451 672
rect -383 638 -371 672
rect -463 632 -371 638
rect -185 672 -93 678
rect -185 638 -173 672
rect -105 638 -93 672
rect -185 632 -93 638
rect 93 672 185 678
rect 93 638 105 672
rect 173 638 185 672
rect 93 632 185 638
rect 371 672 463 678
rect 371 638 383 672
rect 451 638 463 672
rect 371 632 463 638
rect 649 672 741 678
rect 649 638 661 672
rect 729 638 741 672
rect 649 632 741 638
rect 927 672 1019 678
rect 927 638 939 672
rect 1007 638 1019 672
rect 927 632 1019 638
rect -1075 588 -1029 600
rect -1075 -588 -1069 588
rect -1035 -588 -1029 588
rect -1075 -600 -1029 -588
rect -917 588 -871 600
rect -917 -588 -911 588
rect -877 -588 -871 588
rect -917 -600 -871 -588
rect -797 588 -751 600
rect -797 -588 -791 588
rect -757 -588 -751 588
rect -797 -600 -751 -588
rect -639 588 -593 600
rect -639 -588 -633 588
rect -599 -588 -593 588
rect -639 -600 -593 -588
rect -519 588 -473 600
rect -519 -588 -513 588
rect -479 -588 -473 588
rect -519 -600 -473 -588
rect -361 588 -315 600
rect -361 -588 -355 588
rect -321 -588 -315 588
rect -361 -600 -315 -588
rect -241 588 -195 600
rect -241 -588 -235 588
rect -201 -588 -195 588
rect -241 -600 -195 -588
rect -83 588 -37 600
rect -83 -588 -77 588
rect -43 -588 -37 588
rect -83 -600 -37 -588
rect 37 588 83 600
rect 37 -588 43 588
rect 77 -588 83 588
rect 37 -600 83 -588
rect 195 588 241 600
rect 195 -588 201 588
rect 235 -588 241 588
rect 195 -600 241 -588
rect 315 588 361 600
rect 315 -588 321 588
rect 355 -588 361 588
rect 315 -600 361 -588
rect 473 588 519 600
rect 473 -588 479 588
rect 513 -588 519 588
rect 473 -600 519 -588
rect 593 588 639 600
rect 593 -588 599 588
rect 633 -588 639 588
rect 593 -600 639 -588
rect 751 588 797 600
rect 751 -588 757 588
rect 791 -588 797 588
rect 751 -600 797 -588
rect 871 588 917 600
rect 871 -588 877 588
rect 911 -588 917 588
rect 871 -600 917 -588
rect 1029 588 1075 600
rect 1029 -588 1035 588
rect 1069 -588 1075 588
rect 1029 -600 1075 -588
rect -1019 -638 -927 -632
rect -1019 -672 -1007 -638
rect -939 -672 -927 -638
rect -1019 -678 -927 -672
rect -741 -638 -649 -632
rect -741 -672 -729 -638
rect -661 -672 -649 -638
rect -741 -678 -649 -672
rect -463 -638 -371 -632
rect -463 -672 -451 -638
rect -383 -672 -371 -638
rect -463 -678 -371 -672
rect -185 -638 -93 -632
rect -185 -672 -173 -638
rect -105 -672 -93 -638
rect -185 -678 -93 -672
rect 93 -638 185 -632
rect 93 -672 105 -638
rect 173 -672 185 -638
rect 93 -678 185 -672
rect 371 -638 463 -632
rect 371 -672 383 -638
rect 451 -672 463 -638
rect 371 -678 463 -672
rect 649 -638 741 -632
rect 649 -672 661 -638
rect 729 -672 741 -638
rect 649 -678 741 -672
rect 927 -638 1019 -632
rect 927 -672 939 -638
rect 1007 -672 1019 -638
rect 927 -678 1019 -672
<< properties >>
string FIXED_BBOX -1186 -793 1186 793
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 6 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
