**.subckt tb_dac_cell2_dc
V1 net1 GND 3.3
V2 net2 GND 3
V3 net3 GND 0.7
V4 net6 net7 0
V5 net5 net4 0
R1 net4 GND 200 m=1
R2 net7 GND 200 m=1
R4 net8 GND 150k m=1
x1 net1 net8 GND net2 net3 net6 net5 dac_cell2
**** begin user architecture code


.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.param mc_pr_switch=0
*** ANALYSIS TO DO

.dc V2 0.1 3.3 0.001
.save i(V4) i(V5)

.control
set wr_vecnames
set wr_singlescale

run
******** results filename  ************ nodes to write
wrdata $DEV_PATH/res/dac_cell1_dc.res i(V4) i(V5)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  dac_cell2.sym # of pins=7
* sym_path: /opt/uniccass/dev/dac_cell2/tb/dac_cell2.sym
* sch_path: /opt/uniccass/dev/dac_cell2/tb/dac_cell2.sch
.subckt dac_cell2  vsup iref vgnd vsw vbias iout_n iout
*.iopin vsup
*.iopin vgnd
*.iopin iref
*.iopin vsw
*.iopin iout
*.iopin iout_n
*.iopin vbias
XM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 net1 iref net2 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 iout vsw net1 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 iout_n vbias net1 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XR1 net3 vsup vgnd sky130_fd_pr__res_iso_pw W=6.5 L=26.5 mult=1 m=1
XR2 net2 net3 vgnd sky130_fd_pr__res_iso_pw W=6.5 L=26.5 mult=1 m=1
XR3 net3 net2 vgnd sky130_fd_pr__res_iso_pw W=6.5 L=26.5 mult=1 m=1
XR4 vsup net3 vgnd sky130_fd_pr__res_iso_pw W=6.5 L=26.5 mult=1 m=1
.ends

.GLOBAL GND
** flattened .save nodes
.save i(V4) i(V5)
.end
