magic
tech sky130A
magscale 1 2
timestamp 1695288709
<< metal1 >>
rect 0 164000 4000 168000
rect 44000 164000 48000 168000
rect 88000 164000 92000 168000
rect 132000 164000 136000 168000
rect 0 0 4000 4000
rect 44000 0 48000 4000
rect 88000 0 92000 4000
rect 132000 0 136000 4000
use dac  dac_0
timestamp 1695199131
transform 1 0 119831 0 1 144764
box -95 -1536 3512 14414
<< labels >>
rlabel metal1 0 164000 4000 168000 1 bit3
rlabel metal1 44000 164000 48000 168000 1 bit2
rlabel metal1 88000 164000 92000 168000 1 bit1
rlabel metal1 132000 164000 136000 168000 1 bit0
rlabel metal1 0 0 4000 4000 1 power
rlabel metal1 44000 0 48000 4000 1 ground
rlabel metal1 88000 0 92000 4000 1 outsig
rlabel metal1 132000 0 136000 4000 1 vsw
<< end >>
