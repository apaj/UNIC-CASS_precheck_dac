* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p69_RV3JGD a_n69_1300# a_n69_n1732# a_n199_n1862#
X0 a_n69_1300# a_n69_n1732# a_n199_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#2 a_n100_n197# a_100_n100# w_n358_n397#
+ a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n358_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGR8VM a_n100_n497# a_100_n400# w_n358_n697#
+ a_n158_n400#
X0 a_100_n400# a_n100_n497# a_n158_n400# w_n358_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt dac_cell3 vsup iref vsw iout iout_n vbias vgnd
XXR1 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69_RV3JGD
XXR2 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69_RV3JGD
XXR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69_RV3JGD
XXR4 vsup parR vgnd sky130_fd_pr__res_xhigh_po_0p69_RV3JGD
XXM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#2
XXM2 iref sourceM3M4 vsup sourceM2 sky130_fd_pr__pfet_g5v0d10v5_FGR8VM
XXM3 vsw iout vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGR8VM
XXM4 vbias iout_n vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGR8VM
.ends

.subckt sky130_fd_pr__res_high_po_5p73_6QQPRG a_n573_125# a_n573_n557# a_n703_n687#
X0 a_n573_125# a_n573_n557# a_n703_n687# sky130_fd_pr__res_high_po_5p73 l=1.25
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_MS44J6 a_n69_n6232# a_n69_5800# a_n199_n6362#
X0 a_n69_5800# a_n69_n6232# a_n199_n6362# sky130_fd_pr__res_xhigh_po_0p69 l=58
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0 a_n100_n197# a_100_n100# w_n358_n397#
+ a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n358_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt dac_cell1 vsup iref vsw iout iout_n vbias vgnd
XXR1 parR sourceM2 vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXR2 parR sourceM2 vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXR4 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69_MS44J6
XXM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0
XXM2 iref sourceM3M4 vsup sourceM2 sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0
XXM3 vsw iout vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0
XXM4 vbias iout_n vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#0
.ends

.subckt sky130_fd_pr__res_xhigh_po_2p85_5DPYAB a_n415_n687# a_n285_125# a_n285_n557#
X0 a_n285_125# a_n285_n557# a_n415_n687# sky130_fd_pr__res_xhigh_po_2p85 l=1.25
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_PZAK34 a_n165_n982# a_n35_n852# a_n35_420#
X0 a_n35_420# a_n35_n852# a_n165_n982# sky130_fd_pr__res_xhigh_po_0p35 l=4.2
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_5CVACY a_n199_n1162# a_n69_600# a_n69_n1032#
X0 a_n69_600# a_n69_n1032# a_n199_n1162# sky130_fd_pr__res_xhigh_po_0p69 l=6
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y a_50_n500# a_n242_n722# a_n108_n500# a_n50_n588#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n242_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NQCFE9 a_189_n500# a_89_n588# a_31_n500# a_n189_n588#
+ a_n381_n722# a_n89_n500# a_n247_n500#
X0 a_189_n500# a_89_n588# a_31_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
X1 a_n89_n500# a_n189_n588# a_n247_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CJGAEC a_189_n500# a_89_n588# a_31_n500# a_n189_n588#
+ a_n381_n722# a_n89_n500# a_n247_n500#
X0 a_189_n500# a_89_n588# a_31_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
X1 a_n89_n500# a_n189_n588# a_n247_n500# a_n381_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2MGL8M a_367_n688# a_89_n688# a_31_n600# a_n189_n688#
+ a_n1023_n688# a_645_n688# a_n467_n688# a_923_n688# a_n745_n688# a_n89_n600# a_n367_n600#
+ a_n645_n600# a_n1081_n600# a_n247_n600# a_n923_n600# a_n525_n600# a_n803_n600# a_309_n600#
+ a_587_n600# a_189_n600# a_865_n600# a_467_n600# a_n1215_n822# a_745_n600# a_1023_n600#
X0 a_n367_n600# a_n467_n688# a_n525_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X1 a_467_n600# a_367_n688# a_309_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X2 a_189_n600# a_89_n688# a_31_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X3 a_n645_n600# a_n745_n688# a_n803_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X4 a_745_n600# a_645_n688# a_587_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X5 a_n89_n600# a_n189_n688# a_n247_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X6 a_n923_n600# a_n1023_n688# a_n1081_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
X7 a_1023_n600# a_923_n688# a_865_n600# a_n1215_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_X3UTN5 a_170_n700# a_n50_n797# a_50_n700# a_n228_n700#
+ w_n586_n997# a_n108_n700# a_n386_n700# a_228_n797# a_n328_n797# a_328_n700#
X0 a_328_n700# a_228_n797# a_170_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X1 a_50_n700# a_n50_n797# a_n108_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X2 a_n228_n700# a_n328_n797# a_n386_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AE43MT a_170_n700# a_n50_n797# a_50_n700# a_n228_n700#
+ w_n586_n997# a_n108_n700# a_n386_n700# a_228_n797# a_n328_n797# a_328_n700#
X0 a_328_n700# a_228_n797# a_170_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X1 a_50_n700# a_n50_n797# a_n108_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
X2 a_n228_n700# a_n328_n797# a_n386_n700# w_n586_n997# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CNRWF7 a_1579_n1300# a_n803_n1300# a_n1757_n1300#
+ a_n2035_n1300# a_1301_n1300# a_n645_n1300# a_1143_n1300# a_n2413_n1397# a_n2691_n1397#
+ a_n1637_n1300# a_n2193_n1300# w_n2949_n1597# a_189_n1300# a_n525_n1300# a_2591_n1397#
+ a_2313_n1397# a_923_n1397# a_2533_n1300# a_1023_n1300# a_n1479_n1300# a_n367_n1300#
+ a_n1201_n1300# a_n1857_n1397# a_n2135_n1397# a_n745_n1397# a_2691_n1300# a_2413_n1300#
+ a_n89_n1300# a_n1359_n1300# a_n247_n1300# a_645_n1397# a_2255_n1300# a_1977_n1300#
+ a_865_n1300# a_2035_n1397# a_1757_n1397# a_n2749_n1300# a_n1579_n1397# a_n1301_n1397#
+ a_2135_n1300# a_1857_n1300# a_745_n1300# a_n467_n1397# a_n1081_n1300# a_n2313_n1300#
+ a_n2591_n1300# a_89_n1397# a_587_n1300# a_309_n1300# a_1479_n1397# a_367_n1397#
+ a_1699_n1300# a_31_n1300# a_n923_n1300# a_1201_n1397# a_1421_n1300# a_n1915_n1300#
+ a_n2471_n1300# a_467_n1300# a_n189_n1397# a_n1023_n1397#
X0 a_1857_n1300# a_1757_n1397# a_1699_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X1 a_2691_n1300# a_2591_n1397# a_2533_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X2 a_n923_n1300# a_n1023_n1397# a_n1081_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X3 a_745_n1300# a_645_n1397# a_587_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X4 a_n2035_n1300# a_n2135_n1397# a_n2193_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X5 a_1579_n1300# a_1479_n1397# a_1421_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X6 a_467_n1300# a_367_n1397# a_309_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X7 a_n645_n1300# a_n745_n1397# a_n803_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X8 a_n2591_n1300# a_n2691_n1397# a_n2749_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X9 a_n1757_n1300# a_n1857_n1397# a_n1915_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X10 a_n367_n1300# a_n467_n1397# a_n525_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X11 a_1301_n1300# a_1201_n1397# a_1143_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X12 a_2413_n1300# a_2313_n1397# a_2255_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X13 a_n1479_n1300# a_n1579_n1397# a_n1637_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X14 a_n89_n1300# a_n189_n1397# a_n247_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X15 a_2135_n1300# a_2035_n1397# a_1977_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X16 a_189_n1300# a_89_n1397# a_31_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X17 a_n1201_n1300# a_n1301_n1397# a_n1359_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X18 a_1023_n1300# a_923_n1397# a_865_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
X19 a_n2313_n1300# a_n2413_n1397# a_n2471_n1300# w_n2949_n1597# sky130_fd_pr__pfet_g5v0d10v5 ad=3.77 pd=26.6 as=3.77 ps=26.6 w=13 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_C5B489 c1_n1050_n1400# m3_n1150_n1500#
X0 c1_n1050_n1400# m3_n1150_n1500# sky130_fd_pr__cap_mim_m3_1 l=14 w=10
.ends

.subckt miel21_opamp inPos inNeg outSingle power ground
XXR1 ground m1_n1838_8400# bias sky130_fd_pr__res_xhigh_po_0p69_5CVACY
XXR2 ground m1_n1838_8400# m1_360_8394# sky130_fd_pr__res_xhigh_po_0p69_5CVACY
XXR3 ground m1_360_8394# power sky130_fd_pr__res_xhigh_po_0p69_5CVACY
XXM1 d1 ground nsources inPos sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM2 d2 ground nsources inNeg sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM3 bias bias ground bias ground bias ground sky130_fd_pr__nfet_g5v0d10v5_NQCFE9
XXM4 nsources bias ground bias ground nsources ground sky130_fd_pr__nfet_g5v0d10v5_CJGAEC
XXM5 bias bias ground bias bias bias bias bias bias outSingle outSingle outSingle
+ ground ground outSingle ground ground ground ground outSingle ground outSingle ground
+ outSingle outSingle sky130_fd_pr__nfet_g5v0d10v5_2MGL8M
XXM6 power d1 d1 d1 power power power d1 d1 d1 sky130_fd_pr__pfet_g5v0d10v5_X3UTN5
XXM7 power d1 d2 d2 power power power d1 d1 d2 sky130_fd_pr__pfet_g5v0d10v5_AE43MT
XXM8 outSingle power outSingle outSingle outSingle outSingle power d2 d2 power power
+ power outSingle power d2 d2 d2 power outSingle outSingle outSingle outSingle d2
+ d2 d2 outSingle outSingle outSingle power power d2 power power power d2 d2 power
+ d2 d2 outSingle outSingle outSingle d2 power outSingle outSingle d2 power power
+ d2 d2 power power outSingle d2 power power power outSingle d2 d2 sky130_fd_pr__pfet_g5v0d10v5_CNRWF7
XXC1 outSingle d2 sky130_fd_pr__cap_mim_m3_1_C5B489
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_C4MSH5 a_n69_630# a_n69_n1062# a_n199_n1192#
X0 a_n69_630# a_n69_n1062# a_n199_n1192# sky130_fd_pr__res_xhigh_po_0p69 l=6.3
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGUWVM a_n100_n197# a_100_n100# w_n358_n397#
+ a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n358_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FG5HVM a_n100_n897# a_100_n800# a_n158_n800#
+ w_n358_n1097#
X0 a_100_n800# a_n100_n897# a_n158_n800# w_n358_n1097# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=2.32 ps=16.6 w=8 l=1
.ends

.subckt dac_cell4 vsup iref vsw iout iout_n vbias vgnd
XXR1 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69_C4MSH5
XXR2 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69_C4MSH5
XXR3 vsup parR vgnd sky130_fd_pr__res_xhigh_po_0p69_C4MSH5
XXR4 vsup parR vgnd sky130_fd_pr__res_xhigh_po_0p69_C4MSH5
XXM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5_FGUWVM
XXM2 iref sourceM3M4 sourceM2 vsup sky130_fd_pr__pfet_g5v0d10v5_FG5HVM
XXM3 vsw iout sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5_FG5HVM
XXM4 vbias iout_n sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5_FG5HVM
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_XZX24Q a_n199_n3262# a_n69_n3132# a_n69_2700#
X0 a_n69_2700# a_n69_n3132# a_n199_n3262# sky130_fd_pr__res_xhigh_po_0p69 l=27
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#1 a_n100_n197# a_100_n100# w_n358_n397#
+ a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n358_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGK6VM a_n100_n297# a_100_n200# w_n358_n497#
+ a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n358_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt dac_cell2 vsup iref vsw iout iout_n vbias vgnd
XXR1 vgnd parR sourceM2 sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR2 vgnd parR sourceM2 sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR3 vgnd parR vsup sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXR4 vgnd parR vsup sky130_fd_pr__res_xhigh_po_0p69_XZX24Q
XXM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#1
XXM2 iref sourceM3M4 vsup sourceM2 sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
XXM3 vsw iout vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
XXM4 vbias iout_n vsup sourceM3M4 sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
.ends

.subckt dac_top_cell in1 in2 in3 in4 vbias07 vgnd vsup out vbias18
Xdac_cell3_0 vsup in_iref in3 vgnd dac_cell4_0/iout_n vbias07 vgnd dac_cell3
Xsky130_fd_pr__res_high_po_5p73_6QQPRG_1 in_iref m1_n10096_n18392# vgnd sky130_fd_pr__res_high_po_5p73_6QQPRG
Xsky130_fd_pr__res_high_po_5p73_6QQPRG_0 in_iref m1_n10096_n18392# vgnd sky130_fd_pr__res_high_po_5p73_6QQPRG
Xdac_cell1_0 vsup in_iref in1 vgnd dac_cell4_0/iout_n vbias07 vgnd dac_cell1
Xsky130_fd_pr__res_high_po_5p73_6QQPRG_2 vgnd m1_n10096_n18392# vgnd sky130_fd_pr__res_high_po_5p73_6QQPRG
XXR1 vgnd m1_n10096_n18392# vgnd sky130_fd_pr__res_high_po_5p73_6QQPRG
XXR2 vgnd op_amp_in m1_8170_n12070# sky130_fd_pr__res_xhigh_po_2p85_5DPYAB
XXR3 vgnd m1_15440_5366# op_amp_in sky130_fd_pr__res_xhigh_po_0p35_PZAK34
Xmiel21_opamp_0 op_amp_in vbias18 out vsup vgnd miel21_opamp
Xdac_cell4_0 vsup in_iref in4 vgnd dac_cell4_0/iout_n vbias07 vgnd dac_cell4
Xdac_cell2_0 vsup in_iref in2 vgnd dac_cell4_0/iout_n vbias07 vgnd dac_cell2
Xsky130_fd_pr__res_xhigh_po_2p85_5DPYAB_0 vgnd dac_cell4_0/iout_n m1_8170_n12070#
+ sky130_fd_pr__res_xhigh_po_2p85_5DPYAB
Xsky130_fd_pr__res_xhigh_po_2p85_5DPYAB_1 vgnd op_amp_in m1_8170_n12070# sky130_fd_pr__res_xhigh_po_2p85_5DPYAB
Xsky130_fd_pr__res_xhigh_po_2p85_5DPYAB_2 vgnd dac_cell4_0/iout_n m1_8170_n12070#
+ sky130_fd_pr__res_xhigh_po_2p85_5DPYAB
Xsky130_fd_pr__res_xhigh_po_0p35_PZAK34_0 vgnd m1_15440_5366# out sky130_fd_pr__res_xhigh_po_0p35_PZAK34
Xsky130_fd_pr__res_xhigh_po_0p35_PZAK34_1 vgnd m1_15440_5366# op_amp_in sky130_fd_pr__res_xhigh_po_0p35_PZAK34
Xsky130_fd_pr__res_xhigh_po_0p35_PZAK34_2 vgnd m1_15440_5366# out sky130_fd_pr__res_xhigh_po_0p35_PZAK34
.ends

.subckt user_analog_proj_example dac_top_cell_0/vsup dac_top_cell_0/out dac_top_cell_0/in4
+ dac_top_cell_0/in3 dac_top_cell_0/in2 dac_top_cell_0/in1 dac_top_cell_0/vbias07
+ dac_top_cell_0/vbias18 VSUBS
Xdac_top_cell_0 dac_top_cell_0/in1 dac_top_cell_0/in2 dac_top_cell_0/in3 dac_top_cell_0/in4
+ dac_top_cell_0/vbias07 VSUBS dac_top_cell_0/vsup dac_top_cell_0/out dac_top_cell_0/vbias18
+ dac_top_cell
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xuser_analog_proj_example_0 io_analog[7] io_analog[3] io_analog[4] io_analog[2] io_analog[1]
+ io_analog[0] io_analog[6] io_analog[5] vssa1 user_analog_proj_example
.ends

