
**.subckt tb_dac_cell
V1 net1 GND 3.3
V2 net2 GND 3
V3 net3 GND 0.7
V4 net6 net7 0
V5 net5 net4 0
R1 net4 GND 200 m=1
R2 net7 GND 200 m=1
x1 net1 GND net8 net5 net6 net2 net3 dac_cell1
R4 net8 GND 300k m=1
**** begin user architecture code


.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.param mc_pr_switch=0
*** ANALYSIS TO DO

.dc V2 0.1 3.3 0.001
.save i(V4) i(V5)

.control
set wr_vecnames
set wr_singlescale

run
******** results filename  ************ nodes to write
wrdata postlayout_dc.res i(V4) i(V5)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  dac_cell.sym # of pins=7
* sym_path: /home/dder/dac_cell/dac_fourth_cell/tb/dac_cell.sym
* sch_path: /home/dder/dac_cell/dac_fourth_cell/tb/dac_cell.sch

*.option scale=5000u

.subckt dac_cell1 vsup vgnd iref iout iout_n vsw vbias
X0 vsup m1_n66_3062# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=440
X1 vsup m1_n66_3062# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=440
X2 m1_704_2192# m1_n66_3062# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=440
X3 m1_704_2192# m1_n66_3062# vgnd sky130_fd_pr__res_xhigh_po_0p69 l=440
X4 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=278400 pd=12384 as=0 ps=0 w=200 l=200
X5 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X6 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X7 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X8 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X9 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X10 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X11 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X12 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X13 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X14 m1_510_694# vsw iout vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=11600 ps=516 w=200 l=200
X15 m1_704_2192# iref m1_510_694# vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X16 m1_510_694# vbias iout_n vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=11600 ps=516 w=200 l=200
X17 vsup iref iref vsup sky130_fd_pr__pfet_g5v0d10v5 ad=11600 pd=516 as=11600 ps=516 w=200 l=200
X18 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
X19 vgnd vgnd vgnd vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=200
.ends

.GLOBAL GND
** flattened .save nodes
.save i(V4) i(V5)
.end
