magic
tech sky130A
magscale 1 2
timestamp 1698216219
<< locali >>
rect -3804 2478 -3582 2570
rect -3804 396 -3740 2478
rect -3644 396 -3582 2478
rect -3804 328 -3582 396
rect -3176 2462 -2954 2562
rect -3176 380 -3118 2462
rect -3022 380 -2954 2462
rect -3176 320 -2954 380
rect -2564 2474 -2342 2562
rect -2564 392 -2510 2474
rect -2414 392 -2342 2474
rect -2564 320 -2342 392
rect -1958 2462 -1736 2554
rect -1958 380 -1890 2462
rect -1794 380 -1736 2462
rect -1958 312 -1736 380
rect -990 852 -814 1830
rect -990 614 -974 852
rect -830 614 -814 852
rect -990 -100 -814 614
rect -4572 -172 -4360 -120
rect -4572 -2714 -4532 -172
rect -4422 -2714 -4360 -172
rect -1186 -160 -814 -100
rect -3776 -410 -3554 -322
rect -3776 -2492 -3714 -410
rect -3618 -2492 -3554 -410
rect -3776 -2564 -3554 -2492
rect -3176 -410 -2954 -318
rect -3176 -2492 -3122 -410
rect -3026 -2492 -2954 -410
rect -3176 -2560 -2954 -2492
rect -2584 -434 -2362 -322
rect -2584 -2516 -2526 -434
rect -2430 -2516 -2362 -434
rect -2584 -2564 -2362 -2516
rect -1984 -414 -1762 -326
rect -1984 -2496 -1930 -414
rect -1834 -2496 -1762 -414
rect -1984 -2568 -1762 -2496
rect -4572 -2766 -4360 -2714
rect -1186 -2702 -1130 -160
rect -1020 -1298 -814 -160
rect -534 862 -358 1832
rect -534 860 -134 862
rect -534 836 -6 860
rect -534 610 -408 836
rect -22 610 -6 836
rect -534 588 -6 610
rect -534 294 424 588
rect -534 218 -118 294
rect -534 -30 -458 218
rect -158 -30 -118 218
rect -534 -260 -118 -30
rect -52 174 26 202
rect -52 -84 -38 174
rect 8 -84 26 174
rect -52 -88 26 -84
rect 240 178 318 208
rect 240 -80 258 178
rect 304 -80 318 178
rect 240 -88 318 -80
rect -54 -168 318 -88
rect -534 -1296 -358 -260
rect -276 -264 -118 -260
rect -1020 -2702 -974 -1298
rect -1186 -2746 -974 -2702
<< viali >>
rect -3740 396 -3644 2478
rect -3118 380 -3022 2462
rect -2510 392 -2414 2474
rect -1890 380 -1794 2462
rect -974 614 -830 852
rect -4532 -2714 -4422 -172
rect -3714 -2492 -3618 -410
rect -3122 -2492 -3026 -410
rect -2526 -2516 -2430 -434
rect -1930 -2496 -1834 -414
rect -1130 -2702 -1020 -160
rect -408 610 -22 836
rect -458 -30 -158 218
rect -38 -84 8 174
rect 258 -80 304 178
<< metal1 >>
rect -3772 2478 -3614 2534
rect -4058 214 -3888 2438
rect -3772 396 -3740 2478
rect -3644 396 -3614 2478
rect -3144 2462 -2986 2514
rect -3772 372 -3614 396
rect -3470 214 -3300 2422
rect -3144 380 -3118 2462
rect -3022 380 -2986 2462
rect -2534 2474 -2376 2510
rect -3144 352 -2986 380
rect -2870 214 -2700 2422
rect -2534 392 -2510 2474
rect -2414 392 -2376 2474
rect -1926 2462 -1768 2518
rect -2534 348 -2376 392
rect -2270 214 -2100 2426
rect -1926 380 -1890 2462
rect -1794 380 -1768 2462
rect -1926 356 -1768 380
rect -1678 214 -1508 2414
rect -990 852 -812 868
rect -990 614 -974 852
rect -830 614 -812 852
rect -990 592 -812 614
rect -754 512 -582 1748
rect -438 836 10 856
rect -438 610 -408 836
rect -22 610 10 836
rect -438 588 10 610
rect 86 512 186 756
rect -754 340 654 512
rect -476 218 -138 234
rect -4874 210 -598 214
rect -4874 -10 -586 210
rect -4580 -172 -4356 -116
rect -4580 -2714 -4532 -172
rect -4422 -2666 -4356 -172
rect -4058 -2420 -3888 -10
rect -3748 -410 -3590 -374
rect -3748 -2492 -3714 -410
rect -3618 -2492 -3590 -410
rect -3470 -2436 -3300 -10
rect -3156 -410 -2998 -382
rect -3748 -2536 -3590 -2492
rect -3156 -2492 -3122 -410
rect -3026 -2492 -2998 -410
rect -2870 -2436 -2700 -10
rect -2548 -434 -2390 -390
rect -3156 -2544 -2998 -2492
rect -2548 -2516 -2526 -434
rect -2430 -2516 -2390 -434
rect -2270 -2432 -2100 -10
rect -1954 -414 -1796 -378
rect -2548 -2552 -2390 -2516
rect -1954 -2496 -1930 -414
rect -1834 -2496 -1796 -414
rect -1678 -2444 -1508 -10
rect -1194 -160 -970 -108
rect -1954 -2540 -1796 -2496
rect -1194 -2666 -1130 -160
rect -4422 -2702 -1130 -2666
rect -1020 -2452 -970 -160
rect -754 -1184 -586 -10
rect -476 -30 -458 218
rect -158 -30 -138 218
rect -476 -44 -138 -30
rect -52 174 26 202
rect -52 -84 -38 174
rect 8 -84 26 174
rect 86 -28 186 340
rect 240 178 318 208
rect -52 -88 26 -84
rect 240 -80 258 178
rect 304 -80 318 178
rect 240 -88 318 -80
rect -54 -168 318 -88
rect -52 -1752 316 -168
rect -52 -2014 -36 -1752
rect 290 -2014 316 -1752
rect -52 -2028 316 -2014
rect -1020 -2702 -972 -2452
rect -4422 -2714 -972 -2702
rect -4580 -2770 -972 -2714
rect -4578 -2846 -972 -2770
<< via1 >>
rect -3740 396 -3644 2478
rect -3118 380 -3022 2462
rect -2510 392 -2414 2474
rect -1890 380 -1794 2462
rect -974 614 -830 852
rect -408 610 -22 836
rect -3714 -2492 -3618 -410
rect -3122 -2492 -3026 -410
rect -2526 -2516 -2430 -434
rect -1930 -2496 -1834 -414
rect -1130 -1600 -1020 -160
rect -458 -30 -158 218
rect -36 -2014 290 -1752
<< metal2 >>
rect -4892 2478 -1000 2614
rect -4892 396 -3740 2478
rect -3644 2474 -1000 2478
rect -3644 2462 -2510 2474
rect -3644 396 -3118 2462
rect -4892 380 -3118 396
rect -3022 392 -2510 2462
rect -2414 2462 -1000 2474
rect -2414 392 -1890 2462
rect -3022 380 -1890 392
rect -1794 864 -1000 2462
rect -1794 852 12 864
rect -1794 614 -974 852
rect -830 836 12 852
rect -830 614 -408 836
rect -1794 610 -408 614
rect -22 610 12 836
rect -1794 588 12 610
rect -1794 380 -1000 588
rect -4892 320 -1000 380
rect -1174 232 -1000 320
rect -1174 218 -136 232
rect -1174 -30 -458 218
rect -158 -30 -136 218
rect -1174 -44 -136 -30
rect -1174 -160 -1000 -44
rect -4858 -410 -1424 -344
rect -4858 -2492 -3714 -410
rect -3618 -2492 -3122 -410
rect -3026 -414 -1424 -410
rect -3026 -434 -1930 -414
rect -3026 -2492 -2526 -434
rect -4858 -2516 -2526 -2492
rect -2430 -2496 -1930 -434
rect -1834 -1730 -1424 -414
rect -1174 -1600 -1130 -160
rect -1020 -1600 -1000 -160
rect -1174 -1624 -1000 -1600
rect -1834 -1752 312 -1730
rect -1834 -2014 -36 -1752
rect 290 -2014 312 -1752
rect -1834 -2034 312 -2014
rect -1834 -2496 -1424 -2034
rect -2430 -2516 -1424 -2496
rect -4858 -2638 -1424 -2516
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  sky130_fd_pr__diode_pd2nw_05v5_K4SERG_0
timestamp 1698167064
transform 1 0 139 0 1 25
box -321 -321 321 321
use sky130_fd_pr__diode_pd2nw_11v0_PWJNKD  sky130_fd_pr__diode_pd2nw_11v0_PWJNKD_0
timestamp 1697634299
transform 1 0 -2772 0 1 -1448
box -1670 -1378 1670 1378
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0
timestamp 1698167064
transform 1 0 131 0 1 711
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_11v0_2UARL4  sky130_fd_pr__diode_pw2nd_11v0_2UARL4_0
timestamp 1697634299
transform 1 0 -2762 0 1 1438
box -1504 -1172 1504 1172
use sky130_fd_pr__res_high_po_0p35_JFN4DV  sky130_fd_pr__res_high_po_0p35_JFN4DV_0
timestamp 1697634299
transform 1 0 -673 0 1 266
box -201 -1598 201 1598
<< labels >>
rlabel metal2 -4840 368 -4648 2548 1 vgnd
port 2 n
rlabel metal1 452 368 638 494 1 gate
port 3 n
rlabel metal1 -4862 16 -4670 208 1 pad
port 1 n
rlabel metal2 -4828 -2572 -4636 -392 1 vsup
port 0 n
<< end >>
