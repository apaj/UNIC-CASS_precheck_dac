magic
tech sky130A
magscale 1 2
timestamp 1697955996
<< pwell >>
rect -235 -1898 235 1898
<< psubdiff >>
rect -199 1828 -103 1862
rect 103 1828 199 1862
rect -199 1766 -165 1828
rect 165 1766 199 1828
rect -199 -1828 -165 -1766
rect 165 -1828 199 -1766
rect -199 -1862 -103 -1828
rect 103 -1862 199 -1828
<< psubdiffcont >>
rect -103 1828 103 1862
rect -199 -1766 -165 1766
rect 165 -1766 199 1766
rect -103 -1862 103 -1828
<< xpolycontact >>
rect -69 1300 69 1732
rect -69 -1732 69 -1300
<< xpolyres >>
rect -69 -1300 69 1300
<< locali >>
rect -199 1828 -103 1862
rect 103 1828 199 1862
rect -199 1766 -165 1828
rect 165 1766 199 1828
rect -199 -1828 -165 -1766
rect 165 -1828 199 -1766
rect -199 -1862 -103 -1828
rect 103 -1862 199 -1828
<< viali >>
rect -53 1317 53 1714
rect -53 -1714 53 -1317
<< metal1 >>
rect -59 1714 59 1726
rect -59 1317 -53 1714
rect 53 1317 59 1714
rect -59 1305 59 1317
rect -59 -1317 59 -1305
rect -59 -1714 -53 -1317
rect 53 -1714 59 -1317
rect -59 -1726 59 -1714
<< res0p69 >>
rect -71 -1302 71 1302
<< properties >>
string FIXED_BBOX -182 -1845 182 1845
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 13.0 m 1 nx 1 wmin 0.690 lmin 0.50 rho 2000 val 38.226k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
