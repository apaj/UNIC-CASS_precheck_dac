magic
tech sky130A
magscale 1 2
timestamp 1697617627
<< viali >>
rect 892 3814 932 4022
rect 908 3324 948 3532
rect 892 2820 932 3028
rect -3490 2534 -3270 2754
rect 906 2312 946 2520
rect -2592 1078 -2322 1112
rect -1674 962 -1528 1108
rect -508 962 -328 1122
rect -1326 472 -1008 506
rect -1328 -148 -1036 -110
rect -162 -160 138 -124
rect -1790 -804 -1666 -634
<< metal1 >>
rect 878 4022 968 4050
rect -2662 3808 -2224 3990
rect -4210 3804 -2224 3808
rect -4310 3780 -2224 3804
rect -4704 3578 -2224 3780
rect -4310 3532 -2224 3578
rect -4310 1494 -3974 3532
rect -2662 3368 -2224 3532
rect -2672 2780 -2238 2998
rect -3526 2754 -2238 2780
rect -3526 2534 -3490 2754
rect -3270 2534 -2238 2754
rect -3526 2516 -2238 2534
rect -2672 2338 -2238 2516
rect 378 2344 802 3990
rect 878 3814 892 4022
rect 932 3814 968 4022
rect 878 3532 968 3814
rect 878 3324 908 3532
rect 948 3324 968 3532
rect 878 3028 968 3324
rect 878 2820 892 3028
rect 932 2820 968 3028
rect 878 2520 968 2820
rect 878 2320 906 2520
rect 852 2312 906 2320
rect 946 2312 968 2520
rect 852 2098 968 2312
rect -2544 1900 -1092 1906
rect -2544 1774 -1090 1900
rect 852 1898 1052 2098
rect -2544 1540 -2350 1774
rect -4310 1484 -3236 1494
rect -2042 1486 -1876 1774
rect -1278 1530 -1090 1774
rect -4310 1310 -2570 1484
rect -2346 1384 -1876 1486
rect -2346 1312 -1874 1384
rect -3866 1308 -2570 1310
rect -3866 516 -3548 1308
rect -2624 1124 -2312 1136
rect -2628 1112 -2312 1124
rect -2628 1078 -2592 1112
rect -2322 1078 -2312 1112
rect -2628 1060 -2312 1078
rect -2628 516 -2322 1060
rect -2066 914 -1874 1312
rect -1718 1108 -1298 1156
rect -1718 962 -1674 1108
rect -1528 962 -1298 1108
rect -1718 926 -1298 962
rect -1080 1122 -292 1158
rect -1080 962 -508 1122
rect -328 962 -292 1122
rect -1080 928 -292 962
rect -1600 922 -1298 926
rect -2066 714 -1866 914
rect -1350 516 -990 542
rect -3868 506 -990 516
rect -3868 472 -1326 506
rect -1008 472 -990 506
rect -3868 440 -990 472
rect -3868 400 -1066 440
rect -3868 398 -2516 400
rect -3866 396 -3548 398
rect -1350 -84 -1066 400
rect -1350 -110 146 -84
rect -1350 -148 -1328 -110
rect -1036 -124 146 -110
rect -1036 -148 -162 -124
rect -1350 -160 -162 -148
rect 138 -160 146 -124
rect -1350 -166 146 -160
rect -1348 -170 146 -166
rect -1314 -172 146 -170
rect -176 -174 146 -172
rect -1864 -634 -1304 -514
rect -1864 -804 -1790 -634
rect -1666 -804 -1304 -634
rect -596 -652 -126 -528
rect -872 -694 -662 -690
rect -1864 -912 -1304 -804
rect -1074 -898 -660 -694
rect -596 -822 -580 -652
rect -456 -822 -126 -652
rect -596 -840 -126 -822
rect -1268 -1720 -1094 -1178
rect -872 -1564 -662 -898
rect 94 -904 508 -700
rect -872 -1702 -652 -1564
rect -104 -1684 70 -1182
rect -1286 -1918 -1090 -1720
rect -1286 -2118 -1084 -1918
rect -852 -2072 -652 -1702
rect -106 -1800 70 -1684
rect 294 -1728 504 -904
rect -106 -2000 94 -1800
rect 296 -1970 502 -1728
<< via1 >>
rect -3490 2534 -3270 2754
rect -1674 962 -1528 1108
rect -508 962 -328 1122
rect -1790 -804 -1666 -634
rect -580 -822 -456 -652
<< metal2 >>
rect -3562 2754 -3216 2794
rect -3562 2534 -3490 2754
rect -3270 2534 -3216 2754
rect -3562 2510 -3216 2534
rect -3558 2140 -3222 2510
rect -3558 1974 -1494 2140
rect -1738 1168 -1494 1974
rect -1738 1108 -1492 1168
rect -1738 962 -1674 1108
rect -1528 962 -1492 1108
rect -1738 916 -1492 962
rect -570 1122 -296 1150
rect -570 962 -508 1122
rect -328 962 -296 1122
rect -1738 910 -1494 916
rect -570 250 -296 962
rect -726 246 -296 250
rect -1848 72 -296 246
rect -1842 -634 -1602 72
rect -1842 -804 -1790 -634
rect -1666 -804 -1602 -634
rect -1842 -832 -1602 -804
rect -1836 -838 -1602 -832
rect -602 -652 -414 72
rect -602 -822 -580 -652
rect -456 -822 -414 -652
rect -602 -840 -414 -822
rect -602 -846 -426 -840
use sky130_fd_pr__pfet_g5v0d10v5_FGUWVM#2  XM1
timestamp 1697388883
transform 1 0 -2458 0 1 1397
box -358 -397 358 397
use sky130_fd_pr__pfet_g5v0d10v5_FGR8VM  XM2
timestamp 1697388883
transform 1 0 -1184 0 1 1087
box -358 -697 358 697
use sky130_fd_pr__pfet_g5v0d10v5_FGR8VM  XM3
timestamp 1697388883
transform 1 0 -1184 0 1 -733
box -358 -697 358 697
use sky130_fd_pr__pfet_g5v0d10v5_FGR8VM  XM4
timestamp 1697388883
transform 1 0 -18 0 1 -743
box -358 -697 358 697
use sky130_fd_pr__res_xhigh_po_0p69_RV3JGD  XR1
timestamp 1697388883
transform 0 -1 -918 1 0 2415
box -235 -1898 235 1898
use sky130_fd_pr__res_xhigh_po_0p69_RV3JGD  XR2
timestamp 1697388883
transform 0 -1 -934 1 0 2925
box -235 -1898 235 1898
use sky130_fd_pr__res_xhigh_po_0p69_RV3JGD  XR3
timestamp 1697388883
transform 0 1 -918 -1 0 3425
box -235 -1898 235 1898
use sky130_fd_pr__res_xhigh_po_0p69_RV3JGD  XR4
timestamp 1697388883
transform 0 -1 -934 1 0 3915
box -235 -1898 235 1898
<< labels >>
flabel metal1 -4704 3578 -4504 3778 0 FreeSans 128 0 0 0 vsup
port 0 nsew
flabel metal1 852 1898 1052 2098 0 FreeSans 128 0 0 0 vgnd
port 1 nsew
flabel metal1 -2066 714 -1866 914 0 FreeSans 128 0 0 0 iref
port 2 nsew
flabel metal1 -1284 -2118 -1084 -1918 0 FreeSans 128 0 0 0 vsw
port 3 nsew
flabel metal1 -852 -2072 -652 -1872 0 FreeSans 128 0 0 0 iout
port 4 nsew
flabel metal1 -106 -2000 94 -1800 0 FreeSans 128 0 0 0 vbias
port 6 nsew
flabel metal1 296 -1970 496 -1770 0 FreeSans 128 0 0 0 iout_n
port 5 nsew
rlabel metal2 -2798 2000 -2144 2110 1 sourceM2
rlabel metal2 -932 106 -438 224 1 sourceM3M4
rlabel metal1 530 2850 616 3466 1 parR
<< end >>
