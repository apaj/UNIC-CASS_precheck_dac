magic
tech sky130A
magscale 1 2
timestamp 1697955996
<< pwell >>
rect -451 -723 451 723
<< psubdiff >>
rect -415 653 -319 687
rect 319 653 415 687
rect -415 591 -381 653
rect 381 591 415 653
rect -415 -653 -381 -591
rect 381 -653 415 -591
rect -415 -687 -319 -653
rect 319 -687 415 -653
<< psubdiffcont >>
rect -319 653 319 687
rect -415 -591 -381 591
rect 381 -591 415 591
rect -319 -687 319 -653
<< xpolycontact >>
rect -285 125 285 557
rect -285 -557 285 -125
<< xpolyres >>
rect -285 -125 285 125
<< locali >>
rect -415 653 -319 687
rect 319 653 415 687
rect -415 591 -381 653
rect 381 591 415 653
rect -415 -653 -381 -591
rect 381 -653 415 -591
rect -415 -687 -319 -653
rect 319 -687 415 -653
<< viali >>
rect -269 142 269 539
rect -269 -539 269 -142
<< metal1 >>
rect -281 539 281 545
rect -281 142 -269 539
rect 269 142 281 539
rect -281 136 281 142
rect -281 -142 281 -136
rect -281 -539 -269 -142
rect 269 -539 281 -142
rect -281 -545 281 -539
<< res2p85 >>
rect -287 -127 287 127
<< properties >>
string FIXED_BBOX -398 -670 398 670
string gencell sky130_fd_pr__res_xhigh_po_2p85
string library sky130
string parameters w 2.850 l 1.25 m 1 nx 1 wmin 2.850 lmin 0.50 rho 2000 val 1.009k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 2.850 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
