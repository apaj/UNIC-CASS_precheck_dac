magic
tech sky130A
magscale 1 2
timestamp 1698012353
<< nwell >>
rect -586 -997 586 997
<< mvpmos >>
rect -328 -700 -228 700
rect -50 -700 50 700
rect 228 -700 328 700
<< mvpdiff >>
rect -386 688 -328 700
rect -386 -688 -374 688
rect -340 -688 -328 688
rect -386 -700 -328 -688
rect -228 688 -170 700
rect -228 -688 -216 688
rect -182 -688 -170 688
rect -228 -700 -170 -688
rect -108 688 -50 700
rect -108 -688 -96 688
rect -62 -688 -50 688
rect -108 -700 -50 -688
rect 50 688 108 700
rect 50 -688 62 688
rect 96 -688 108 688
rect 50 -700 108 -688
rect 170 688 228 700
rect 170 -688 182 688
rect 216 -688 228 688
rect 170 -700 228 -688
rect 328 688 386 700
rect 328 -688 340 688
rect 374 -688 386 688
rect 328 -700 386 -688
<< mvpdiffc >>
rect -374 -688 -340 688
rect -216 -688 -182 688
rect -96 -688 -62 688
rect 62 -688 96 688
rect 182 -688 216 688
rect 340 -688 374 688
<< mvnsubdiff >>
rect -520 919 520 931
rect -520 885 -412 919
rect 412 885 520 919
rect -520 873 520 885
rect -520 823 -462 873
rect -520 -823 -508 823
rect -474 -823 -462 823
rect 462 823 520 873
rect -520 -873 -462 -823
rect 462 -823 474 823
rect 508 -823 520 823
rect 462 -873 520 -823
rect -520 -885 520 -873
rect -520 -919 -412 -885
rect 412 -919 520 -885
rect -520 -931 520 -919
<< mvnsubdiffcont >>
rect -412 885 412 919
rect -508 -823 -474 823
rect 474 -823 508 823
rect -412 -919 412 -885
<< poly >>
rect -328 781 -228 797
rect -328 747 -312 781
rect -244 747 -228 781
rect -328 700 -228 747
rect -50 781 50 797
rect -50 747 -34 781
rect 34 747 50 781
rect -50 700 50 747
rect 228 781 328 797
rect 228 747 244 781
rect 312 747 328 781
rect 228 700 328 747
rect -328 -747 -228 -700
rect -328 -781 -312 -747
rect -244 -781 -228 -747
rect -328 -797 -228 -781
rect -50 -747 50 -700
rect -50 -781 -34 -747
rect 34 -781 50 -747
rect -50 -797 50 -781
rect 228 -747 328 -700
rect 228 -781 244 -747
rect 312 -781 328 -747
rect 228 -797 328 -781
<< polycont >>
rect -312 747 -244 781
rect -34 747 34 781
rect 244 747 312 781
rect -312 -781 -244 -747
rect -34 -781 34 -747
rect 244 -781 312 -747
<< locali >>
rect -508 885 -412 919
rect 412 885 508 919
rect -508 823 -474 885
rect 474 823 508 885
rect -328 747 -312 781
rect -244 747 -228 781
rect -50 747 -34 781
rect 34 747 50 781
rect 228 747 244 781
rect 312 747 328 781
rect -374 688 -340 704
rect -374 -704 -340 -688
rect -216 688 -182 704
rect -216 -704 -182 -688
rect -96 688 -62 704
rect -96 -704 -62 -688
rect 62 688 96 704
rect 62 -704 96 -688
rect 182 688 216 704
rect 182 -704 216 -688
rect 340 688 374 704
rect 340 -704 374 -688
rect -328 -781 -312 -747
rect -244 -781 -228 -747
rect -50 -781 -34 -747
rect 34 -781 50 -747
rect 228 -781 244 -747
rect 312 -781 328 -747
rect -508 -885 -474 -823
rect 474 -885 508 -823
rect -508 -919 -412 -885
rect 412 -919 508 -885
<< viali >>
rect -312 747 -244 781
rect -34 747 34 781
rect 244 747 312 781
rect -374 -688 -340 688
rect -216 -688 -182 688
rect -96 -688 -62 688
rect 62 -688 96 688
rect 182 -688 216 688
rect 340 -688 374 688
rect -312 -781 -244 -747
rect -34 -781 34 -747
rect 244 -781 312 -747
<< metal1 >>
rect -324 781 -232 787
rect -324 747 -312 781
rect -244 747 -232 781
rect -324 741 -232 747
rect -46 781 46 787
rect -46 747 -34 781
rect 34 747 46 781
rect -46 741 46 747
rect 232 781 324 787
rect 232 747 244 781
rect 312 747 324 781
rect 232 741 324 747
rect -380 688 -334 700
rect -380 -688 -374 688
rect -340 -688 -334 688
rect -380 -700 -334 -688
rect -222 688 -176 700
rect -222 -688 -216 688
rect -182 -688 -176 688
rect -222 -700 -176 -688
rect -102 688 -56 700
rect -102 -688 -96 688
rect -62 -688 -56 688
rect -102 -700 -56 -688
rect 56 688 102 700
rect 56 -688 62 688
rect 96 -688 102 688
rect 56 -700 102 -688
rect 176 688 222 700
rect 176 -688 182 688
rect 216 -688 222 688
rect 176 -700 222 -688
rect 334 688 380 700
rect 334 -688 340 688
rect 374 -688 380 688
rect 334 -700 380 -688
rect -324 -747 -232 -741
rect -324 -781 -312 -747
rect -244 -781 -232 -747
rect -324 -787 -232 -781
rect -46 -747 46 -741
rect -46 -781 -34 -747
rect 34 -781 46 -747
rect -46 -787 46 -781
rect 232 -747 324 -741
rect 232 -781 244 -747
rect 312 -781 324 -747
rect 232 -787 324 -781
<< properties >>
string FIXED_BBOX -491 -902 491 902
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 7 l 0.50 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
