magic
tech sky130A
magscale 1 2
timestamp 1697533315
<< pwell >>
rect -831 -858 831 858
<< mvnmos >>
rect -603 -600 -503 600
rect -445 -600 -345 600
rect -287 -600 -187 600
rect -129 -600 -29 600
rect 29 -600 129 600
rect 187 -600 287 600
rect 345 -600 445 600
rect 503 -600 603 600
<< mvndiff >>
rect -661 588 -603 600
rect -661 -588 -649 588
rect -615 -588 -603 588
rect -661 -600 -603 -588
rect -503 588 -445 600
rect -503 -588 -491 588
rect -457 -588 -445 588
rect -503 -600 -445 -588
rect -345 588 -287 600
rect -345 -588 -333 588
rect -299 -588 -287 588
rect -345 -600 -287 -588
rect -187 588 -129 600
rect -187 -588 -175 588
rect -141 -588 -129 588
rect -187 -600 -129 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 129 588 187 600
rect 129 -588 141 588
rect 175 -588 187 588
rect 129 -600 187 -588
rect 287 588 345 600
rect 287 -588 299 588
rect 333 -588 345 588
rect 287 -600 345 -588
rect 445 588 503 600
rect 445 -588 457 588
rect 491 -588 503 588
rect 445 -600 503 -588
rect 603 588 661 600
rect 603 -588 615 588
rect 649 -588 661 588
rect 603 -600 661 -588
<< mvndiffc >>
rect -649 -588 -615 588
rect -491 -588 -457 588
rect -333 -588 -299 588
rect -175 -588 -141 588
rect -17 -588 17 588
rect 141 -588 175 588
rect 299 -588 333 588
rect 457 -588 491 588
rect 615 -588 649 588
<< mvpsubdiff >>
rect -795 810 795 822
rect -795 776 -687 810
rect 687 776 795 810
rect -795 764 795 776
rect -795 714 -737 764
rect -795 -714 -783 714
rect -749 -714 -737 714
rect 737 714 795 764
rect -795 -764 -737 -714
rect 737 -714 749 714
rect 783 -714 795 714
rect 737 -764 795 -714
rect -795 -776 795 -764
rect -795 -810 -687 -776
rect 687 -810 795 -776
rect -795 -822 795 -810
<< mvpsubdiffcont >>
rect -687 776 687 810
rect -783 -714 -749 714
rect 749 -714 783 714
rect -687 -810 687 -776
<< poly >>
rect -603 672 -503 688
rect -603 638 -587 672
rect -519 638 -503 672
rect -603 600 -503 638
rect -445 672 -345 688
rect -445 638 -429 672
rect -361 638 -345 672
rect -445 600 -345 638
rect -287 672 -187 688
rect -287 638 -271 672
rect -203 638 -187 672
rect -287 600 -187 638
rect -129 672 -29 688
rect -129 638 -113 672
rect -45 638 -29 672
rect -129 600 -29 638
rect 29 672 129 688
rect 29 638 45 672
rect 113 638 129 672
rect 29 600 129 638
rect 187 672 287 688
rect 187 638 203 672
rect 271 638 287 672
rect 187 600 287 638
rect 345 672 445 688
rect 345 638 361 672
rect 429 638 445 672
rect 345 600 445 638
rect 503 672 603 688
rect 503 638 519 672
rect 587 638 603 672
rect 503 600 603 638
rect -603 -638 -503 -600
rect -603 -672 -587 -638
rect -519 -672 -503 -638
rect -603 -688 -503 -672
rect -445 -638 -345 -600
rect -445 -672 -429 -638
rect -361 -672 -345 -638
rect -445 -688 -345 -672
rect -287 -638 -187 -600
rect -287 -672 -271 -638
rect -203 -672 -187 -638
rect -287 -688 -187 -672
rect -129 -638 -29 -600
rect -129 -672 -113 -638
rect -45 -672 -29 -638
rect -129 -688 -29 -672
rect 29 -638 129 -600
rect 29 -672 45 -638
rect 113 -672 129 -638
rect 29 -688 129 -672
rect 187 -638 287 -600
rect 187 -672 203 -638
rect 271 -672 287 -638
rect 187 -688 287 -672
rect 345 -638 445 -600
rect 345 -672 361 -638
rect 429 -672 445 -638
rect 345 -688 445 -672
rect 503 -638 603 -600
rect 503 -672 519 -638
rect 587 -672 603 -638
rect 503 -688 603 -672
<< polycont >>
rect -587 638 -519 672
rect -429 638 -361 672
rect -271 638 -203 672
rect -113 638 -45 672
rect 45 638 113 672
rect 203 638 271 672
rect 361 638 429 672
rect 519 638 587 672
rect -587 -672 -519 -638
rect -429 -672 -361 -638
rect -271 -672 -203 -638
rect -113 -672 -45 -638
rect 45 -672 113 -638
rect 203 -672 271 -638
rect 361 -672 429 -638
rect 519 -672 587 -638
<< locali >>
rect -783 776 -687 810
rect 687 776 783 810
rect -783 714 -749 776
rect 749 714 783 776
rect -603 638 -587 672
rect -519 638 -503 672
rect -445 638 -429 672
rect -361 638 -345 672
rect -287 638 -271 672
rect -203 638 -187 672
rect -129 638 -113 672
rect -45 638 -29 672
rect 29 638 45 672
rect 113 638 129 672
rect 187 638 203 672
rect 271 638 287 672
rect 345 638 361 672
rect 429 638 445 672
rect 503 638 519 672
rect 587 638 603 672
rect -649 588 -615 604
rect -649 -604 -615 -588
rect -491 588 -457 604
rect -491 -604 -457 -588
rect -333 588 -299 604
rect -333 -604 -299 -588
rect -175 588 -141 604
rect -175 -604 -141 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 141 588 175 604
rect 141 -604 175 -588
rect 299 588 333 604
rect 299 -604 333 -588
rect 457 588 491 604
rect 457 -604 491 -588
rect 615 588 649 604
rect 615 -604 649 -588
rect -603 -672 -587 -638
rect -519 -672 -503 -638
rect -445 -672 -429 -638
rect -361 -672 -345 -638
rect -287 -672 -271 -638
rect -203 -672 -187 -638
rect -129 -672 -113 -638
rect -45 -672 -29 -638
rect 29 -672 45 -638
rect 113 -672 129 -638
rect 187 -672 203 -638
rect 271 -672 287 -638
rect 345 -672 361 -638
rect 429 -672 445 -638
rect 503 -672 519 -638
rect 587 -672 603 -638
rect -783 -776 -749 -714
rect 749 -776 783 -714
rect -783 -810 -687 -776
rect 687 -810 783 -776
<< viali >>
rect -587 638 -519 672
rect -429 638 -361 672
rect -271 638 -203 672
rect -113 638 -45 672
rect 45 638 113 672
rect 203 638 271 672
rect 361 638 429 672
rect 519 638 587 672
rect -649 -588 -615 588
rect -491 -588 -457 588
rect -333 -588 -299 588
rect -175 -588 -141 588
rect -17 -588 17 588
rect 141 -588 175 588
rect 299 -588 333 588
rect 457 -588 491 588
rect 615 -588 649 588
rect -587 -672 -519 -638
rect -429 -672 -361 -638
rect -271 -672 -203 -638
rect -113 -672 -45 -638
rect 45 -672 113 -638
rect 203 -672 271 -638
rect 361 -672 429 -638
rect 519 -672 587 -638
<< metal1 >>
rect -599 672 -507 678
rect -599 638 -587 672
rect -519 638 -507 672
rect -599 632 -507 638
rect -441 672 -349 678
rect -441 638 -429 672
rect -361 638 -349 672
rect -441 632 -349 638
rect -283 672 -191 678
rect -283 638 -271 672
rect -203 638 -191 672
rect -283 632 -191 638
rect -125 672 -33 678
rect -125 638 -113 672
rect -45 638 -33 672
rect -125 632 -33 638
rect 33 672 125 678
rect 33 638 45 672
rect 113 638 125 672
rect 33 632 125 638
rect 191 672 283 678
rect 191 638 203 672
rect 271 638 283 672
rect 191 632 283 638
rect 349 672 441 678
rect 349 638 361 672
rect 429 638 441 672
rect 349 632 441 638
rect 507 672 599 678
rect 507 638 519 672
rect 587 638 599 672
rect 507 632 599 638
rect -655 588 -609 600
rect -655 -588 -649 588
rect -615 -588 -609 588
rect -655 -600 -609 -588
rect -497 588 -451 600
rect -497 -588 -491 588
rect -457 -588 -451 588
rect -497 -600 -451 -588
rect -339 588 -293 600
rect -339 -588 -333 588
rect -299 -588 -293 588
rect -339 -600 -293 -588
rect -181 588 -135 600
rect -181 -588 -175 588
rect -141 -588 -135 588
rect -181 -600 -135 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 135 588 181 600
rect 135 -588 141 588
rect 175 -588 181 588
rect 135 -600 181 -588
rect 293 588 339 600
rect 293 -588 299 588
rect 333 -588 339 588
rect 293 -600 339 -588
rect 451 588 497 600
rect 451 -588 457 588
rect 491 -588 497 588
rect 451 -600 497 -588
rect 609 588 655 600
rect 609 -588 615 588
rect 649 -588 655 588
rect 609 -600 655 -588
rect -599 -638 -507 -632
rect -599 -672 -587 -638
rect -519 -672 -507 -638
rect -599 -678 -507 -672
rect -441 -638 -349 -632
rect -441 -672 -429 -638
rect -361 -672 -349 -638
rect -441 -678 -349 -672
rect -283 -638 -191 -632
rect -283 -672 -271 -638
rect -203 -672 -191 -638
rect -283 -678 -191 -672
rect -125 -638 -33 -632
rect -125 -672 -113 -638
rect -45 -672 -33 -638
rect -125 -678 -33 -672
rect 33 -638 125 -632
rect 33 -672 45 -638
rect 113 -672 125 -638
rect 33 -678 125 -672
rect 191 -638 283 -632
rect 191 -672 203 -638
rect 271 -672 283 -638
rect 191 -678 283 -672
rect 349 -638 441 -632
rect 349 -672 361 -638
rect 429 -672 441 -638
rect 349 -678 441 -672
rect 507 -638 599 -632
rect 507 -672 519 -638
rect 587 -672 599 -638
rect 507 -678 599 -672
<< properties >>
string FIXED_BBOX -766 -793 766 793
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 6.0 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
