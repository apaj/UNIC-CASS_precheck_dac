magic
tech sky130A
magscale 1 2
timestamp 1697533315
<< metal3 >>
rect -1150 1472 1149 1500
rect -1150 -1472 1065 1472
rect 1129 -1472 1149 1472
rect -1150 -1500 1149 -1472
<< via3 >>
rect 1065 -1472 1129 1472
<< mimcap >>
rect -1050 1360 950 1400
rect -1050 -1360 -1010 1360
rect 910 -1360 950 1360
rect -1050 -1400 950 -1360
<< mimcapcontact >>
rect -1010 -1360 910 1360
<< metal4 >>
rect 1049 1472 1145 1488
rect -1011 1360 911 1361
rect -1011 -1360 -1010 1360
rect 910 -1360 911 1360
rect -1011 -1361 911 -1360
rect 1049 -1472 1065 1472
rect 1129 -1472 1145 1472
rect 1049 -1488 1145 -1472
<< properties >>
string FIXED_BBOX -1150 -1500 1050 1500
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 14.0 val 289.12 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
