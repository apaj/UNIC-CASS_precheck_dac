* SPICE3 file created from dac_cell2.ext - technology: sky130A

.option scale=5000u

*.subckt dac_cell2 vsup vgnd iref vsw iout iout_n vbias
*.iopin vsup
*.iopin vgnd
*.iopin iref
*.iopin vsw
*.iopin iout
*.iopin iout_n
*.iopin vbias
X0 net2 net3 vgnd sky130_fd_pr__res_xhigh_po_0p69 l=5400
X1 net2 net3 vgnd sky130_fd_pr__res_xhigh_po_0p69 l=5400
X2 net3 vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=5400
X3 net3 vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 l=5400
X4 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 ad=11600 pd=516 as=11600 ps=516 w=200 l=200
X5 net1 iref net2 vsup sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=400 l=200
X6 iout vsw net1 vsup sky130_fd_pr__pfet_g5v0d10v5 ad=23200 pd=916 as=0 ps=0 w=400 l=200
X7 iout_n vbias net1 vsup sky130_fd_pr__pfet_g5v0d10v5 ad=23200 pd=916 as=0 ps=0 w=400 l=200
*.ends
** flattened .save nodes
*.end
