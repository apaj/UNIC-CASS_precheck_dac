magic
tech sky130A
magscale 1 2
timestamp 1697955996
<< nwell >>
rect 730 6170 1290 8170
<< psubdiff >>
rect -1110 2820 -800 2850
rect -1110 2680 -1080 2820
rect -830 2680 -800 2820
rect -1110 2650 -800 2680
<< psubdiffcont >>
rect -1080 2680 -830 2820
<< viali >>
rect -648 8756 -428 8796
rect -642 8630 -422 8670
rect -1952 8142 -1918 8292
rect -406 7126 -368 7362
rect -218 7126 -180 7362
rect 760 7190 804 7446
rect 1206 7198 1250 7454
rect -672 6038 -462 6078
rect -118 6030 92 6070
rect 648 6022 858 6062
rect -962 5758 -920 5958
rect -1666 5582 -1628 5728
rect -664 3510 -626 3678
rect -1100 2820 -810 2840
rect -1100 2680 -1080 2820
rect -1080 2680 -830 2820
rect -830 2680 -810 2820
rect -1100 2660 -810 2680
<< metal1 >>
rect -1922 9824 -1718 10290
rect -1922 9798 -1570 9824
rect -1922 9692 -1704 9798
rect -1600 9692 -1570 9798
rect -1922 9674 -1570 9692
rect -1922 9024 -1718 9674
rect 1374 9100 6792 9172
rect -1922 8882 -834 9024
rect -668 8796 -410 8814
rect -668 8758 -648 8796
rect -2140 8756 -648 8758
rect -428 8756 -410 8796
rect -2140 8670 -410 8756
rect -2140 8644 -642 8670
rect -2140 8310 -1972 8644
rect -668 8630 -642 8644
rect -422 8630 -410 8670
rect -668 8608 -410 8630
rect -1838 8400 -844 8538
rect -2140 8292 -1908 8310
rect -2140 8142 -1952 8292
rect -1918 8142 -1908 8292
rect -2140 8128 -1908 8142
rect -2140 6230 -1972 8128
rect -1826 7974 -1674 8400
rect 360 8394 782 9030
rect 1342 8976 1410 8986
rect 1342 8716 1350 8976
rect 1402 8716 1410 8976
rect 1342 8706 1410 8716
rect 1610 8974 1680 8984
rect 1610 8714 1620 8974
rect 1672 8714 1680 8974
rect 1610 8708 1680 8714
rect 1892 8974 1960 8990
rect 1892 8714 1900 8974
rect 1952 8714 1960 8974
rect 1892 8710 1960 8714
rect 2164 8974 2232 8982
rect 2164 8714 2174 8974
rect 2226 8714 2232 8974
rect 2164 8702 2232 8714
rect 2444 8974 2512 8982
rect 2444 8714 2454 8974
rect 2506 8714 2512 8974
rect 2444 8702 2512 8714
rect 2724 8974 2792 8986
rect 2724 8714 2732 8974
rect 2784 8714 2792 8974
rect 2724 8706 2792 8714
rect 3000 8974 3068 8986
rect 3000 8714 3010 8974
rect 3062 8714 3068 8974
rect 3000 8706 3068 8714
rect 3284 8974 3352 8982
rect 3284 8714 3290 8974
rect 3342 8714 3352 8974
rect 3284 8702 3352 8714
rect 3558 8974 3626 8980
rect 3558 8714 3566 8974
rect 3618 8714 3626 8974
rect 3558 8700 3626 8714
rect 3834 8974 3902 8984
rect 3834 8714 3844 8974
rect 3896 8714 3902 8974
rect 3834 8704 3902 8714
rect 4114 8974 4182 8986
rect 4114 8714 4122 8974
rect 4174 8714 4182 8974
rect 4114 8706 4182 8714
rect 4392 8974 4460 8980
rect 4392 8714 4400 8974
rect 4452 8714 4460 8974
rect 4392 8700 4460 8714
rect 4668 8974 4736 8984
rect 4668 8714 4678 8974
rect 4730 8714 4736 8974
rect 4668 8704 4736 8714
rect 4950 8974 5018 8984
rect 4950 8714 4956 8974
rect 5008 8714 5018 8974
rect 4950 8704 5018 8714
rect 5224 8974 5292 8986
rect 5224 8714 5234 8974
rect 5286 8714 5292 8974
rect 5224 8706 5292 8714
rect 5506 8974 5574 8984
rect 5506 8714 5512 8974
rect 5564 8714 5574 8974
rect 5506 8704 5574 8714
rect 5780 8974 5848 8988
rect 5780 8714 5788 8974
rect 5840 8714 5848 8974
rect 5780 8708 5848 8714
rect 6068 8974 6120 8982
rect 5788 8706 5840 8708
rect 6068 8706 6120 8714
rect 6346 8974 6398 8982
rect 6346 8706 6398 8714
rect 6622 8974 6680 8982
rect 6674 8714 6680 8974
rect 6622 8706 6680 8714
rect 1766 8492 1842 8502
rect 1496 8478 1572 8484
rect 1496 8218 1502 8478
rect 1554 8218 1572 8478
rect 1766 8232 1774 8492
rect 1826 8232 1842 8492
rect 1766 8222 1842 8232
rect 2040 8498 2116 8504
rect 2040 8238 2056 8498
rect 2108 8238 2116 8498
rect 2040 8224 2116 8238
rect 2322 8496 2398 8506
rect 2322 8236 2332 8496
rect 2384 8236 2398 8496
rect 2322 8226 2398 8236
rect 2602 8496 2678 8504
rect 2602 8236 2610 8496
rect 2662 8236 2678 8496
rect 2602 8224 2678 8236
rect 2876 8496 2952 8506
rect 2876 8236 2890 8496
rect 2942 8236 2952 8496
rect 2876 8226 2952 8236
rect 3152 8496 3228 8506
rect 3152 8236 3166 8496
rect 3218 8236 3228 8496
rect 3152 8226 3228 8236
rect 3434 8496 3510 8510
rect 3434 8236 3446 8496
rect 3498 8236 3510 8496
rect 3434 8230 3510 8236
rect 3708 8496 3784 8506
rect 3708 8236 3722 8496
rect 3774 8236 3784 8496
rect 3708 8226 3784 8236
rect 3992 8496 4068 8504
rect 3992 8236 4000 8496
rect 4052 8236 4068 8496
rect 3992 8224 4068 8236
rect 4266 8496 4342 8504
rect 4266 8236 4278 8496
rect 4330 8236 4342 8496
rect 4266 8224 4342 8236
rect 4544 8496 4620 8506
rect 4544 8236 4556 8496
rect 4608 8236 4620 8496
rect 4544 8226 4620 8236
rect 4826 8496 4902 8506
rect 4826 8236 4836 8496
rect 4888 8236 4902 8496
rect 4826 8226 4902 8236
rect 5102 8496 5178 8508
rect 5102 8236 5112 8496
rect 5164 8236 5178 8496
rect 5102 8228 5178 8236
rect 5380 8496 5456 8504
rect 5380 8236 5392 8496
rect 5444 8236 5456 8496
rect 5380 8224 5456 8236
rect 5658 8496 5734 8508
rect 5658 8236 5668 8496
rect 5720 8236 5734 8496
rect 5658 8228 5734 8236
rect 5936 8496 6012 8508
rect 5936 8236 5946 8496
rect 5998 8236 6012 8496
rect 5936 8228 6012 8236
rect 6214 8496 6290 8506
rect 6214 8236 6226 8496
rect 6278 8236 6290 8496
rect 6214 8226 6290 8236
rect 6492 8496 6560 8504
rect 6492 8236 6502 8496
rect 6554 8236 6560 8496
rect 6492 8224 6560 8236
rect 6772 8496 6840 8506
rect 6772 8236 6780 8496
rect 6832 8236 6840 8496
rect 6772 8226 6840 8236
rect 1496 8204 1572 8218
rect -630 8006 -426 8032
rect -630 8004 -536 8006
rect -632 7956 -536 8004
rect -1208 7934 -536 7956
rect -462 7934 -426 8006
rect -1208 7920 -426 7934
rect -162 8000 50 8022
rect -162 7932 -140 8000
rect -62 7952 50 8000
rect -62 7932 622 7952
rect -1208 7916 -550 7920
rect -162 7912 622 7932
rect -1266 7770 -1202 7780
rect -1266 7508 -1258 7770
rect -1206 7508 -1202 7770
rect -1266 7500 -1202 7508
rect -990 7770 -926 7778
rect -990 7508 -982 7770
rect -930 7508 -926 7770
rect -990 7498 -926 7508
rect -708 7770 -644 7780
rect -708 7508 -704 7770
rect -652 7508 -644 7770
rect -708 7500 -644 7508
rect -98 7750 -28 7776
rect -98 7490 -88 7750
rect -36 7490 -28 7750
rect -98 7484 -28 7490
rect 184 7770 254 7776
rect 184 7510 190 7770
rect 242 7510 254 7770
rect 184 7484 254 7510
rect 458 7770 528 7778
rect 458 7510 468 7770
rect 520 7510 528 7770
rect 458 7486 528 7510
rect 468 7484 526 7486
rect 742 7454 1272 7482
rect 742 7446 1206 7454
rect -430 7362 -148 7398
rect -430 7126 -406 7362
rect -368 7126 -218 7362
rect -180 7126 -148 7362
rect 742 7190 760 7446
rect 804 7334 1206 7446
rect 804 7206 972 7334
rect 1122 7206 1206 7334
rect 804 7198 1206 7206
rect 1250 7198 1272 7454
rect 804 7190 1272 7198
rect 742 7184 1272 7190
rect -430 7106 -148 7126
rect -1108 6932 -1040 6946
rect -1108 6670 -1098 6932
rect -1046 6670 -1040 6932
rect -1108 6664 -1040 6670
rect -830 6932 -768 6944
rect -830 6670 -824 6932
rect -772 6670 -768 6932
rect -830 6664 -768 6670
rect -552 6940 -490 6944
rect -552 6934 -488 6940
rect -552 6672 -546 6934
rect -494 6672 -488 6934
rect -552 6664 -488 6672
rect 58 6916 122 6926
rect 58 6656 68 6916
rect 120 6656 122 6916
rect 58 6650 122 6656
rect 342 6916 406 6924
rect 342 6656 346 6916
rect 398 6656 406 6916
rect 342 6648 406 6656
rect 622 6916 686 6926
rect 622 6656 626 6916
rect 678 6656 686 6916
rect 622 6650 686 6656
rect 942 6432 1466 6436
rect 3586 6432 3772 6434
rect -1222 6382 -530 6432
rect -54 6380 638 6430
rect 942 6420 6782 6432
rect 942 6368 962 6420
rect 1026 6402 6782 6420
rect 1026 6386 3632 6402
rect 1026 6368 1050 6386
rect 1392 6382 3632 6386
rect 942 6348 1050 6368
rect 3586 6332 3632 6382
rect 3712 6382 6782 6402
rect 3712 6332 3772 6382
rect 3586 6308 3772 6332
rect -2058 5970 -1974 6230
rect 58 6100 880 6106
rect -980 6094 880 6100
rect -982 6078 880 6094
rect -982 6038 -672 6078
rect -462 6070 880 6078
rect -462 6038 -118 6070
rect -982 6030 -118 6038
rect 92 6062 880 6070
rect 92 6030 648 6062
rect -982 6024 648 6030
rect -1342 5978 -1256 5984
rect -2058 5950 -1770 5970
rect -2058 5868 -1922 5950
rect -1812 5868 -1770 5950
rect -1342 5948 -1336 5978
rect -1494 5922 -1336 5948
rect -1264 5948 -1256 5978
rect -982 5958 -876 6024
rect -682 6022 648 6024
rect 858 6022 880 6062
rect -682 6008 880 6022
rect 58 5996 880 6008
rect 9100 6078 9690 6172
rect -1264 5922 -1090 5948
rect -1494 5900 -1090 5922
rect -2058 5846 -1770 5868
rect -1548 5814 -1476 5820
rect -1682 5732 -1598 5770
rect -1682 5604 -1670 5732
rect -1616 5604 -1598 5732
rect -1682 5582 -1666 5604
rect -1628 5582 -1598 5604
rect -1682 5564 -1598 5582
rect -1548 5554 -1538 5814
rect -1482 5554 -1476 5814
rect -1548 5548 -1476 5554
rect -1274 5814 -1184 5824
rect -1274 5554 -1260 5814
rect -1204 5554 -1184 5814
rect -982 5758 -962 5958
rect -920 5758 -876 5958
rect -982 5752 -876 5758
rect -694 5828 -624 5834
rect -694 5568 -688 5828
rect -630 5568 -624 5828
rect -694 5562 -624 5568
rect -128 5820 -58 5826
rect -128 5560 -122 5820
rect -64 5560 -58 5820
rect -128 5554 -58 5560
rect 458 5806 544 5822
rect -1274 5550 -1184 5554
rect -1260 5548 -1198 5550
rect 458 5546 474 5806
rect 530 5546 544 5806
rect 458 5534 544 5546
rect 744 5806 816 5814
rect 744 5546 752 5806
rect 808 5546 816 5806
rect 744 5538 816 5546
rect 1020 5806 1092 5816
rect 1020 5546 1028 5806
rect 1084 5546 1092 5806
rect 1020 5540 1092 5546
rect 1298 5806 1370 5814
rect 1298 5546 1306 5806
rect 1362 5546 1370 5806
rect 1298 5538 1370 5546
rect 1576 5806 1648 5814
rect 1576 5546 1584 5806
rect 1640 5546 1648 5806
rect 1576 5538 1648 5546
rect 1856 5806 1928 5814
rect 1856 5546 1864 5806
rect 1920 5546 1928 5806
rect 1856 5538 1928 5546
rect 2134 5806 2206 5814
rect 2134 5546 2142 5806
rect 2198 5546 2206 5806
rect 2134 5538 2206 5546
rect 2412 5806 2484 5814
rect 2412 5546 2420 5806
rect 2476 5546 2484 5806
rect 2412 5538 2484 5546
rect 9100 5792 9172 6078
rect 9524 5792 9690 6078
rect 9100 5366 9690 5792
rect -1402 5224 -1314 5246
rect -1402 4964 -1380 5224
rect -1324 4964 -1314 5224
rect -1402 4940 -1314 4964
rect -1120 5224 -1032 5256
rect -1120 4964 -1102 5224
rect -1046 4964 -1032 5224
rect -536 5234 -466 5240
rect -536 4972 -530 5234
rect -472 4972 -466 5234
rect -536 4966 -466 4972
rect 30 5234 100 5240
rect 30 4972 36 5234
rect 94 4972 100 5234
rect 30 4966 100 4972
rect 622 5014 694 5022
rect -1120 4950 -1032 4964
rect -3490 4738 -2778 4856
rect -1484 4788 -1106 4836
rect -624 4828 -540 4830
rect -3490 4444 -3170 4738
rect -2876 4444 -2778 4738
rect -3490 4438 -2778 4444
rect -3488 4436 -3288 4438
rect -1328 4414 -1252 4788
rect -624 4762 -614 4828
rect -544 4762 -540 4828
rect -624 4734 -540 4762
rect -466 4822 -378 4824
rect -466 4778 36 4822
rect -1020 4700 -930 4704
rect -1020 4648 -1008 4700
rect -944 4698 -930 4700
rect -944 4696 -682 4698
rect -466 4696 -378 4778
rect 622 4754 630 5014
rect 688 4754 694 5014
rect 622 4746 694 4754
rect 900 5014 972 5022
rect 900 4754 908 5014
rect 966 4754 972 5014
rect 900 4746 972 4754
rect 1178 5014 1250 5024
rect 1178 4754 1186 5014
rect 1244 4754 1250 5014
rect 1178 4748 1250 4754
rect 1456 5014 1528 5022
rect 1456 4754 1464 5014
rect 1522 4754 1528 5014
rect 1456 4746 1528 4754
rect 1734 5014 1806 5024
rect 1734 4754 1742 5014
rect 1800 4754 1806 5014
rect 1734 4748 1806 4754
rect 2014 5014 2086 5022
rect 2014 4754 2020 5014
rect 2078 4754 2086 5014
rect 2014 4746 2086 4754
rect 2290 5014 2362 5020
rect 2290 4754 2298 5014
rect 2356 4754 2362 5014
rect 2290 4744 2362 4754
rect 2568 5014 2640 5022
rect 2568 4754 2576 5014
rect 2634 4754 2640 5014
rect 2568 4746 2640 4754
rect -944 4672 -378 4696
rect -944 4648 -380 4672
rect -1020 4646 -380 4648
rect -1020 4640 -930 4646
rect -718 4644 -380 4646
rect -126 4512 -20 4678
rect 526 4610 2576 4614
rect 524 4568 2576 4610
rect -2218 4406 -2076 4410
rect -2218 4402 -1556 4406
rect -2218 4396 -1420 4402
rect -2218 4324 -1516 4396
rect -1438 4324 -1420 4396
rect -1328 4372 -100 4414
rect -2218 4312 -1420 4324
rect -2218 3984 -2076 4312
rect -542 4280 -474 4290
rect -542 4020 -536 4280
rect -480 4020 -474 4280
rect -542 4016 -474 4020
rect -266 4286 -198 4290
rect -266 4280 -196 4286
rect -266 4020 -258 4280
rect -202 4020 -196 4280
rect -266 4016 -196 4020
rect -542 4014 -480 4016
rect -258 4014 -196 4016
rect -3488 3980 -2076 3984
rect -3496 3782 -2076 3980
rect -3496 3780 -2190 3782
rect -684 3686 -608 3694
rect -684 3502 -676 3686
rect -616 3502 -608 3686
rect -684 3498 -608 3502
rect -390 3634 -312 3652
rect -390 3374 -376 3634
rect -320 3374 -312 3634
rect -390 3366 -312 3374
rect -108 3636 -30 3652
rect -108 3376 -100 3636
rect -44 3376 -30 3636
rect -108 3366 -30 3376
rect -2332 3098 -2068 3122
rect -2332 2922 -2292 3098
rect -2096 3024 -2068 3098
rect 524 3024 638 4568
rect -2096 2922 638 3024
rect -2332 2892 638 2922
rect -1120 2840 -790 2860
rect -1120 2660 -1100 2840
rect -810 2660 -790 2840
rect -1880 2630 -1628 2648
rect -1120 2640 -790 2660
rect -1880 2468 -1850 2630
rect -1640 2468 -1628 2630
rect -1880 2212 -1628 2468
<< via1 >>
rect -1704 9692 -1600 9798
rect 1350 8716 1402 8976
rect 1620 8714 1672 8974
rect 1900 8714 1952 8974
rect 2174 8714 2226 8974
rect 2454 8714 2506 8974
rect 2732 8714 2784 8974
rect 3010 8714 3062 8974
rect 3290 8714 3342 8974
rect 3566 8714 3618 8974
rect 3844 8714 3896 8974
rect 4122 8714 4174 8974
rect 4400 8714 4452 8974
rect 4678 8714 4730 8974
rect 4956 8714 5008 8974
rect 5234 8714 5286 8974
rect 5512 8714 5564 8974
rect 5788 8714 5840 8974
rect 6068 8714 6120 8974
rect 6346 8714 6398 8974
rect 6622 8714 6674 8974
rect 1502 8218 1554 8478
rect 1774 8232 1826 8492
rect 2056 8238 2108 8498
rect 2332 8236 2384 8496
rect 2610 8236 2662 8496
rect 2890 8236 2942 8496
rect 3166 8236 3218 8496
rect 3446 8236 3498 8496
rect 3722 8236 3774 8496
rect 4000 8236 4052 8496
rect 4278 8236 4330 8496
rect 4556 8236 4608 8496
rect 4836 8236 4888 8496
rect 5112 8236 5164 8496
rect 5392 8236 5444 8496
rect 5668 8236 5720 8496
rect 5946 8236 5998 8496
rect 6226 8236 6278 8496
rect 6502 8236 6554 8496
rect 6780 8236 6832 8496
rect -536 7934 -462 8006
rect -140 7932 -62 8000
rect -1258 7508 -1206 7770
rect -982 7508 -930 7770
rect -704 7508 -652 7770
rect -88 7490 -36 7750
rect 190 7510 242 7770
rect 468 7510 520 7770
rect 972 7206 1122 7334
rect -1804 6366 -1706 6682
rect -1098 6670 -1046 6932
rect -824 6670 -772 6932
rect -546 6672 -494 6934
rect 68 6656 120 6916
rect 346 6656 398 6916
rect 626 6656 678 6916
rect 962 6368 1026 6420
rect 3632 6332 3712 6402
rect -1922 5868 -1812 5950
rect -1336 5922 -1264 5978
rect -1670 5728 -1616 5732
rect -1670 5604 -1666 5728
rect -1666 5604 -1628 5728
rect -1628 5604 -1616 5728
rect -1538 5554 -1482 5814
rect -1260 5554 -1204 5814
rect -688 5568 -630 5828
rect -122 5560 -64 5820
rect 474 5546 530 5806
rect 752 5546 808 5806
rect 1028 5546 1084 5806
rect 1306 5546 1362 5806
rect 1584 5546 1640 5806
rect 1864 5546 1920 5806
rect 2142 5546 2198 5806
rect 2420 5546 2476 5806
rect 9172 5792 9524 6078
rect -1380 4964 -1324 5224
rect -1102 4964 -1046 5224
rect -530 4972 -472 5234
rect 36 4972 94 5234
rect -3170 4444 -2876 4738
rect -614 4762 -544 4828
rect -1008 4648 -944 4700
rect 630 4754 688 5014
rect 908 4754 966 5014
rect 1186 4754 1244 5014
rect 1464 4754 1522 5014
rect 1742 4754 1800 5014
rect 2020 4754 2078 5014
rect 2298 4754 2356 5014
rect 2576 4754 2634 5014
rect -1516 4324 -1438 4396
rect -536 4020 -480 4280
rect -258 4020 -202 4280
rect -676 3678 -616 3686
rect -676 3510 -664 3678
rect -664 3510 -626 3678
rect -626 3510 -616 3678
rect -676 3502 -616 3510
rect -376 3374 -320 3634
rect -100 3376 -44 3636
rect -2292 2922 -2096 3098
rect -1080 2680 -830 2820
rect -1850 2468 -1640 2630
<< metal2 >>
rect 1314 9824 1540 9836
rect -1720 9798 1558 9824
rect -1720 9692 -1704 9798
rect -1600 9692 1558 9798
rect -1720 9674 1558 9692
rect -1420 9554 1558 9674
rect -1420 9548 242 9554
rect -1420 8170 -1292 9548
rect -1420 8044 -1290 8170
rect -1420 7790 -1292 8044
rect -548 8014 -432 8016
rect -548 8006 -52 8014
rect -548 7934 -536 8006
rect -462 8000 -52 8006
rect -462 7934 -140 8000
rect -548 7932 -140 7934
rect -62 7932 -52 8000
rect -548 7926 -52 7932
rect -1420 7770 -636 7790
rect -1420 7508 -1258 7770
rect -1206 7508 -982 7770
rect -930 7508 -704 7770
rect -652 7508 -636 7770
rect -1420 7500 -636 7508
rect -1416 7496 -636 7500
rect -548 6964 -432 7926
rect 98 7788 242 9548
rect -116 7770 540 7788
rect -116 7750 190 7770
rect -116 7490 -88 7750
rect -36 7510 190 7750
rect 242 7510 468 7770
rect 520 7510 540 7770
rect -36 7490 540 7510
rect -116 7478 540 7490
rect 944 7334 1148 9554
rect 1314 9502 1558 9554
rect 1314 9026 1540 9502
rect 1270 8976 6868 9026
rect 1270 8716 1350 8976
rect 1402 8974 6868 8976
rect 1402 8716 1620 8974
rect 1270 8714 1620 8716
rect 1672 8714 1900 8974
rect 1952 8714 2174 8974
rect 2226 8714 2454 8974
rect 2506 8714 2732 8974
rect 2784 8714 3010 8974
rect 3062 8714 3290 8974
rect 3342 8714 3566 8974
rect 3618 8714 3844 8974
rect 3896 8714 4122 8974
rect 4174 8714 4400 8974
rect 4452 8714 4678 8974
rect 4730 8714 4956 8974
rect 5008 8714 5234 8974
rect 5286 8714 5512 8974
rect 5564 8714 5788 8974
rect 5840 8714 6068 8974
rect 6120 8714 6346 8974
rect 6398 8714 6622 8974
rect 6674 8714 6868 8974
rect 1270 8686 6868 8714
rect 1398 8504 7798 8530
rect 1398 8498 8244 8504
rect 1398 8492 2056 8498
rect 1398 8478 1774 8492
rect 1398 8218 1502 8478
rect 1554 8232 1774 8478
rect 1826 8238 2056 8492
rect 2108 8496 8244 8498
rect 2108 8238 2332 8496
rect 1826 8236 2332 8238
rect 2384 8236 2610 8496
rect 2662 8236 2890 8496
rect 2942 8236 3166 8496
rect 3218 8236 3446 8496
rect 3498 8236 3722 8496
rect 3774 8236 4000 8496
rect 4052 8236 4278 8496
rect 4330 8236 4556 8496
rect 4608 8236 4836 8496
rect 4888 8236 5112 8496
rect 5164 8236 5392 8496
rect 5444 8236 5668 8496
rect 5720 8236 5946 8496
rect 5998 8236 6226 8496
rect 6278 8236 6502 8496
rect 6554 8236 6780 8496
rect 6832 8236 8244 8496
rect 1826 8232 8244 8236
rect 1554 8218 8244 8232
rect 1398 8200 8244 8218
rect 1398 8160 8240 8200
rect 944 7206 972 7334
rect 1122 7206 1148 7334
rect 944 7188 1148 7206
rect -1118 6934 -432 6964
rect -1118 6932 -546 6934
rect -1852 6682 -1658 6736
rect -1852 6366 -1804 6682
rect -1706 6366 -1658 6682
rect -1118 6670 -1098 6932
rect -1046 6670 -824 6932
rect -772 6672 -546 6932
rect -494 6672 -432 6934
rect -772 6670 -432 6672
rect -1118 6658 -432 6670
rect 44 6916 690 6934
rect -1852 6348 -1658 6366
rect -2310 6130 -2072 6134
rect -1852 6130 -1656 6348
rect -1102 6146 -1048 6148
rect -2310 6118 -1656 6130
rect -1328 6118 -1048 6146
rect -2310 6040 -1252 6118
rect -3230 4742 -2682 4924
rect -3230 4738 -3146 4742
rect -3230 4444 -3170 4738
rect -3230 4380 -3146 4444
rect -2790 4380 -2682 4742
rect -3230 4188 -2682 4380
rect -2310 3098 -2072 6040
rect -1852 6038 -1252 6040
rect -1816 6036 -1252 6038
rect -1346 5978 -1254 6036
rect -1972 5950 -1770 5978
rect -1972 5868 -1922 5950
rect -1812 5868 -1770 5950
rect -1346 5922 -1336 5978
rect -1264 5922 -1254 5978
rect -1346 5916 -1254 5922
rect -1972 5764 -1770 5868
rect -1560 5814 -1180 5830
rect -1560 5764 -1538 5814
rect -1974 5732 -1538 5764
rect -1974 5604 -1670 5732
rect -1616 5604 -1538 5732
rect -1974 5570 -1538 5604
rect -1974 4282 -1764 5570
rect -1560 5554 -1538 5570
rect -1482 5554 -1260 5814
rect -1204 5554 -1180 5814
rect -1560 5548 -1180 5554
rect -1102 5290 -1048 6118
rect -1422 5224 -1028 5290
rect -856 5236 -724 6658
rect 44 6656 68 6916
rect 120 6656 346 6916
rect 398 6656 626 6916
rect 678 6656 690 6916
rect 44 6646 690 6656
rect 152 6226 320 6646
rect 940 6420 1052 6436
rect 940 6368 962 6420
rect 1026 6368 1052 6420
rect 940 6226 1052 6368
rect 3610 6412 3736 6426
rect 3610 6320 3620 6412
rect 3720 6320 3736 6412
rect 3610 6308 3736 6320
rect 152 6130 1052 6226
rect -694 5828 -624 5834
rect -694 5568 -688 5828
rect -630 5826 -64 5828
rect -630 5820 -58 5826
rect -630 5572 -122 5820
rect -630 5568 -624 5572
rect -694 5562 -624 5568
rect -536 5236 -466 5240
rect -1422 4964 -1380 5224
rect -1324 4964 -1102 5224
rect -1046 4964 -1028 5224
rect -1422 4938 -1028 4964
rect -876 5234 -458 5236
rect -876 4972 -530 5234
rect -472 4974 -458 5234
rect -472 4972 -460 4974
rect -876 4952 -460 4972
rect -624 4828 -534 4838
rect -624 4762 -614 4828
rect -544 4762 -534 4828
rect -1482 4700 -930 4712
rect -1482 4648 -1008 4700
rect -944 4648 -930 4700
rect -1482 4640 -930 4648
rect -1482 4422 -1400 4640
rect -624 4558 -534 4762
rect -364 4648 -228 5572
rect -128 5560 -122 5572
rect -64 5560 -58 5820
rect -128 5554 -58 5560
rect 152 5242 320 6130
rect 7794 6096 8240 8160
rect 7794 6078 9544 6096
rect 7794 5928 9172 6078
rect 32 5240 320 5242
rect 30 5234 320 5240
rect 30 4972 36 5234
rect 94 4980 320 5234
rect 358 5838 466 5842
rect 358 5806 2498 5838
rect 358 5546 474 5806
rect 530 5546 752 5806
rect 808 5546 1028 5806
rect 1084 5546 1306 5806
rect 1362 5546 1584 5806
rect 1640 5546 1864 5806
rect 1920 5546 2142 5806
rect 2198 5546 2420 5806
rect 2476 5546 2498 5806
rect 358 5526 2498 5546
rect 6780 5792 9172 5928
rect 9524 5792 9544 6078
rect 6780 5772 9544 5792
rect 6780 5770 8240 5772
rect 94 4972 242 4980
rect 30 4970 242 4972
rect 30 4966 100 4970
rect -364 4568 214 4648
rect -344 4558 214 4568
rect -920 4546 -534 4558
rect -920 4466 -908 4546
rect -806 4466 -534 4546
rect -920 4454 -534 4466
rect -1522 4396 -1398 4422
rect -1522 4324 -1516 4396
rect -1438 4324 -1398 4396
rect -1522 4320 -1398 4324
rect -542 4282 -194 4296
rect -1974 4280 -194 4282
rect -1974 4022 -536 4280
rect -1974 3714 -1764 4022
rect -542 4020 -536 4022
rect -480 4020 -258 4280
rect -202 4020 -194 4280
rect -542 4012 -194 4020
rect -1974 3688 -604 3714
rect -1978 3686 -604 3688
rect -1978 3502 -676 3686
rect -616 3502 -604 3686
rect -1978 3486 -604 3502
rect -396 3636 -30 3664
rect 78 3636 208 4558
rect 358 4248 466 5526
rect 6780 5260 7110 5770
rect 7628 5260 8240 5770
rect 6780 5078 8240 5260
rect 582 5014 2648 5042
rect 582 4754 630 5014
rect 688 4754 908 5014
rect 966 4754 1186 5014
rect 1244 4754 1464 5014
rect 1522 4754 1742 5014
rect 1800 4754 2020 5014
rect 2078 4754 2298 5014
rect 2356 4754 2576 5014
rect 2634 4754 2648 5014
rect 582 4694 2648 4754
rect 362 3880 458 4248
rect -396 3634 -100 3636
rect -1978 3412 -1762 3486
rect -2310 2922 -2292 3098
rect -2096 2922 -2072 3098
rect -2310 2910 -2072 2922
rect -1974 2840 -1764 3412
rect -396 3374 -376 3634
rect -320 3376 -100 3634
rect -44 3388 210 3636
rect -44 3376 -30 3388
rect -320 3374 -30 3376
rect -396 3350 -30 3374
rect -1120 2840 -790 2860
rect 358 2840 458 3880
rect -1974 2820 458 2840
rect -1974 2680 -1080 2820
rect -830 2680 458 2820
rect -1974 2666 458 2680
rect 2260 4166 2630 4694
rect -1974 2662 436 2666
rect -1974 2630 -1564 2662
rect -1120 2640 -790 2662
rect -1974 2468 -1850 2630
rect -1640 2468 -1564 2630
rect 2260 2548 2632 4166
rect 7794 2548 8240 5078
rect -1974 2462 -1564 2468
rect -1884 2454 -1564 2462
rect 2240 2124 8244 2548
rect 7794 2114 8240 2124
<< via2 >>
rect -3146 4738 -2790 4742
rect -3146 4444 -2876 4738
rect -2876 4444 -2790 4738
rect -3146 4380 -2790 4444
rect 3620 6402 3720 6412
rect 3620 6332 3632 6402
rect 3632 6332 3712 6402
rect 3712 6332 3720 6402
rect 3620 6320 3720 6332
rect -908 4466 -806 4546
rect 7110 5260 7628 5770
<< metal3 >>
rect 3574 6412 3758 6430
rect 3574 6408 3620 6412
rect 3720 6408 3758 6412
rect 3574 6272 3586 6408
rect 3740 6272 3758 6408
rect 3574 6262 3758 6272
rect 6794 5808 7808 5936
rect 6794 5178 6928 5808
rect 7642 5178 7808 5808
rect 6794 5106 7808 5178
rect -3176 4742 -2772 4774
rect -3176 4380 -3146 4742
rect -2790 4560 -2772 4742
rect -2790 4546 -794 4560
rect -2790 4466 -908 4546
rect -806 4466 -794 4546
rect -2790 4454 -794 4466
rect -2790 4380 -2772 4454
rect -3176 4360 -2772 4380
<< via3 >>
rect 3586 6320 3620 6408
rect 3620 6320 3720 6408
rect 3720 6320 3740 6408
rect 3586 6272 3740 6320
rect 6928 5770 7642 5808
rect 6928 5260 7110 5770
rect 7110 5260 7628 5770
rect 7628 5260 7642 5770
rect 6928 5178 7642 5260
<< metal4 >>
rect 3574 6412 3756 6428
rect 3574 6408 5124 6412
rect 3574 6272 3586 6408
rect 3740 6282 5124 6408
rect 3740 6272 5116 6282
rect 3574 6262 5116 6272
rect 3586 6228 5116 6262
rect 5000 5984 5116 6228
rect 6928 5828 7786 5942
rect 6802 5808 7786 5828
rect 6802 5178 6928 5808
rect 7642 5178 7786 5808
rect 6802 5044 7786 5178
rect 4198 3004 4678 4552
rect 6802 3004 7592 5044
rect 4198 2924 7592 3004
rect 4198 2718 7578 2924
rect 4198 2710 4678 2718
use sky130_fd_pr__cap_mim_m3_1_C5B489  XC1
timestamp 1697955996
transform 1 0 3962 0 1 4642
box -1150 -1500 1149 1500
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM1
timestamp 1697955996
transform 1 0 -580 0 1 5364
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM2
timestamp 1697955996
transform 1 0 -14 0 1 5356
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_NQCFE9  XM3
timestamp 1697955996
transform 1 0 -1293 0 1 5364
box -417 -758 417 758
use sky130_fd_pr__nfet_g5v0d10v5_CJGAEC  XM4
timestamp 1697955996
transform 1 0 -289 0 1 3836
box -417 -758 417 758
use sky130_fd_pr__nfet_g5v0d10v5_2MGL8M  XM5
timestamp 1697955996
transform 1 0 1553 0 1 5246
box -1251 -858 1251 858
use sky130_fd_pr__pfet_g5v0d10v5_X3UTN5  XM6
timestamp 1697955996
transform 1 0 -876 0 1 7171
box -586 -997 586 997
use sky130_fd_pr__pfet_g5v0d10v5_AE43MT  XM7
timestamp 1697955996
transform 1 0 294 0 1 7169
box -586 -997 586 997
use sky130_fd_pr__pfet_g5v0d10v5_CNRWF7  XM8
timestamp 1697955996
transform 1 0 4087 0 1 7771
box -2949 -1597 2949 1597
use sky130_fd_pr__res_xhigh_po_0p69_5CVACY  XR1
timestamp 1697955996
transform 1 0 -1751 0 1 7372
box -235 -1198 235 1198
use sky130_fd_pr__res_xhigh_po_0p69_5CVACY  XR2
timestamp 1697955996
transform 0 -1 -240 1 0 8467
box -235 -1198 235 1198
use sky130_fd_pr__res_xhigh_po_0p69_5CVACY  XR3
timestamp 1697955996
transform 0 1 -244 -1 0 8955
box -235 -1198 235 1198
<< labels >>
flabel metal1 -1920 10086 -1720 10286 0 FreeSans 1280 0 0 0 power
port 3 nsew
flabel metal1 -1880 2212 -1680 2412 0 FreeSans 1280 0 0 0 ground
port 4 nsew
flabel metal1 -3488 4436 -3288 4636 0 FreeSans 1280 0 0 0 inPos
port 0 nsew
flabel metal1 -3496 3780 -3296 3980 0 FreeSans 1280 0 0 0 inNeg
port 1 nsew
flabel metal1 9482 5368 9682 5568 0 FreeSans 1280 0 0 0 outSingle
port 2 nsew
rlabel metal2 -1830 6044 -1746 6156 1 bias
rlabel metal2 112 4114 196 4226 1 nsources
rlabel metal2 -828 6062 -744 6174 1 d1
rlabel metal2 184 6050 268 6162 1 d2
<< end >>
