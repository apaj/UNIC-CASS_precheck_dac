magic
tech sky130A
magscale 1 2
timestamp 1628235263
<< pwell >>
rect -673 -5058 673 5058
<< nnmos >>
rect -445 -4800 -345 4800
rect -287 -4800 -187 4800
rect -129 -4800 -29 4800
rect 29 -4800 129 4800
rect 187 -4800 287 4800
rect 345 -4800 445 4800
<< mvndiff >>
rect -503 4788 -445 4800
rect -503 -4788 -491 4788
rect -457 -4788 -445 4788
rect -503 -4800 -445 -4788
rect -345 4788 -287 4800
rect -345 -4788 -333 4788
rect -299 -4788 -287 4788
rect -345 -4800 -287 -4788
rect -187 4788 -129 4800
rect -187 -4788 -175 4788
rect -141 -4788 -129 4788
rect -187 -4800 -129 -4788
rect -29 4788 29 4800
rect -29 -4788 -17 4788
rect 17 -4788 29 4788
rect -29 -4800 29 -4788
rect 129 4788 187 4800
rect 129 -4788 141 4788
rect 175 -4788 187 4788
rect 129 -4800 187 -4788
rect 287 4788 345 4800
rect 287 -4788 299 4788
rect 333 -4788 345 4788
rect 287 -4800 345 -4788
rect 445 4788 503 4800
rect 445 -4788 457 4788
rect 491 -4788 503 4788
rect 445 -4800 503 -4788
<< mvndiffc >>
rect -491 -4788 -457 4788
rect -333 -4788 -299 4788
rect -175 -4788 -141 4788
rect -17 -4788 17 4788
rect 141 -4788 175 4788
rect 299 -4788 333 4788
rect 457 -4788 491 4788
<< mvpsubdiff >>
rect -637 5010 637 5022
rect -637 4976 -529 5010
rect 529 4976 637 5010
rect -637 4964 637 4976
rect -637 4914 -579 4964
rect -637 -4914 -625 4914
rect -591 -4914 -579 4914
rect 579 4914 637 4964
rect -637 -4964 -579 -4914
rect 579 -4914 591 4914
rect 625 -4914 637 4914
rect 579 -4964 637 -4914
rect -637 -4976 637 -4964
rect -637 -5010 -529 -4976
rect 529 -5010 637 -4976
rect -637 -5022 637 -5010
<< mvpsubdiffcont >>
rect -529 4976 529 5010
rect -625 -4914 -591 4914
rect 591 -4914 625 4914
rect -529 -5010 529 -4976
<< poly >>
rect -445 4872 -345 4888
rect -445 4838 -429 4872
rect -361 4838 -345 4872
rect -445 4800 -345 4838
rect -287 4872 -187 4888
rect -287 4838 -271 4872
rect -203 4838 -187 4872
rect -287 4800 -187 4838
rect -129 4872 -29 4888
rect -129 4838 -113 4872
rect -45 4838 -29 4872
rect -129 4800 -29 4838
rect 29 4872 129 4888
rect 29 4838 45 4872
rect 113 4838 129 4872
rect 29 4800 129 4838
rect 187 4872 287 4888
rect 187 4838 203 4872
rect 271 4838 287 4872
rect 187 4800 287 4838
rect 345 4872 445 4888
rect 345 4838 361 4872
rect 429 4838 445 4872
rect 345 4800 445 4838
rect -445 -4838 -345 -4800
rect -445 -4872 -429 -4838
rect -361 -4872 -345 -4838
rect -445 -4888 -345 -4872
rect -287 -4838 -187 -4800
rect -287 -4872 -271 -4838
rect -203 -4872 -187 -4838
rect -287 -4888 -187 -4872
rect -129 -4838 -29 -4800
rect -129 -4872 -113 -4838
rect -45 -4872 -29 -4838
rect -129 -4888 -29 -4872
rect 29 -4838 129 -4800
rect 29 -4872 45 -4838
rect 113 -4872 129 -4838
rect 29 -4888 129 -4872
rect 187 -4838 287 -4800
rect 187 -4872 203 -4838
rect 271 -4872 287 -4838
rect 187 -4888 287 -4872
rect 345 -4838 445 -4800
rect 345 -4872 361 -4838
rect 429 -4872 445 -4838
rect 345 -4888 445 -4872
<< polycont >>
rect -429 4838 -361 4872
rect -271 4838 -203 4872
rect -113 4838 -45 4872
rect 45 4838 113 4872
rect 203 4838 271 4872
rect 361 4838 429 4872
rect -429 -4872 -361 -4838
rect -271 -4872 -203 -4838
rect -113 -4872 -45 -4838
rect 45 -4872 113 -4838
rect 203 -4872 271 -4838
rect 361 -4872 429 -4838
<< locali >>
rect -625 4976 -529 5010
rect 529 4976 625 5010
rect -625 4914 -591 4976
rect 591 4914 625 4976
rect -445 4838 -429 4872
rect -361 4838 -345 4872
rect -287 4838 -271 4872
rect -203 4838 -187 4872
rect -129 4838 -113 4872
rect -45 4838 -29 4872
rect 29 4838 45 4872
rect 113 4838 129 4872
rect 187 4838 203 4872
rect 271 4838 287 4872
rect 345 4838 361 4872
rect 429 4838 445 4872
rect -491 4788 -457 4804
rect -491 -4804 -457 -4788
rect -333 4788 -299 4804
rect -333 -4804 -299 -4788
rect -175 4788 -141 4804
rect -175 -4804 -141 -4788
rect -17 4788 17 4804
rect -17 -4804 17 -4788
rect 141 4788 175 4804
rect 141 -4804 175 -4788
rect 299 4788 333 4804
rect 299 -4804 333 -4788
rect 457 4788 491 4804
rect 457 -4804 491 -4788
rect -445 -4872 -429 -4838
rect -361 -4872 -345 -4838
rect -287 -4872 -271 -4838
rect -203 -4872 -187 -4838
rect -129 -4872 -113 -4838
rect -45 -4872 -29 -4838
rect 29 -4872 45 -4838
rect 113 -4872 129 -4838
rect 187 -4872 203 -4838
rect 271 -4872 287 -4838
rect 345 -4872 361 -4838
rect 429 -4872 445 -4838
rect -625 -4976 -591 -4914
rect 591 -4976 625 -4914
rect -625 -5010 -529 -4976
rect 529 -5010 625 -4976
<< viali >>
rect -429 4838 -361 4872
rect -271 4838 -203 4872
rect -113 4838 -45 4872
rect 45 4838 113 4872
rect 203 4838 271 4872
rect 361 4838 429 4872
rect -491 -4788 -457 4788
rect -333 -4788 -299 4788
rect -175 -4788 -141 4788
rect -17 -4788 17 4788
rect 141 -4788 175 4788
rect 299 -4788 333 4788
rect 457 -4788 491 4788
rect -429 -4872 -361 -4838
rect -271 -4872 -203 -4838
rect -113 -4872 -45 -4838
rect 45 -4872 113 -4838
rect 203 -4872 271 -4838
rect 361 -4872 429 -4838
<< metal1 >>
rect -441 4872 -349 4878
rect -441 4838 -429 4872
rect -361 4838 -349 4872
rect -441 4832 -349 4838
rect -283 4872 -191 4878
rect -283 4838 -271 4872
rect -203 4838 -191 4872
rect -283 4832 -191 4838
rect -125 4872 -33 4878
rect -125 4838 -113 4872
rect -45 4838 -33 4872
rect -125 4832 -33 4838
rect 33 4872 125 4878
rect 33 4838 45 4872
rect 113 4838 125 4872
rect 33 4832 125 4838
rect 191 4872 283 4878
rect 191 4838 203 4872
rect 271 4838 283 4872
rect 191 4832 283 4838
rect 349 4872 441 4878
rect 349 4838 361 4872
rect 429 4838 441 4872
rect 349 4832 441 4838
rect -497 4788 -451 4800
rect -497 -4788 -491 4788
rect -457 -4788 -451 4788
rect -497 -4800 -451 -4788
rect -339 4788 -293 4800
rect -339 -4788 -333 4788
rect -299 -4788 -293 4788
rect -339 -4800 -293 -4788
rect -181 4788 -135 4800
rect -181 -4788 -175 4788
rect -141 -4788 -135 4788
rect -181 -4800 -135 -4788
rect -23 4788 23 4800
rect -23 -4788 -17 4788
rect 17 -4788 23 4788
rect -23 -4800 23 -4788
rect 135 4788 181 4800
rect 135 -4788 141 4788
rect 175 -4788 181 4788
rect 135 -4800 181 -4788
rect 293 4788 339 4800
rect 293 -4788 299 4788
rect 333 -4788 339 4788
rect 293 -4800 339 -4788
rect 451 4788 497 4800
rect 451 -4788 457 4788
rect 491 -4788 497 4788
rect 451 -4800 497 -4788
rect -441 -4838 -349 -4832
rect -441 -4872 -429 -4838
rect -361 -4872 -349 -4838
rect -441 -4878 -349 -4872
rect -283 -4838 -191 -4832
rect -283 -4872 -271 -4838
rect -203 -4872 -191 -4838
rect -283 -4878 -191 -4872
rect -125 -4838 -33 -4832
rect -125 -4872 -113 -4838
rect -45 -4872 -33 -4838
rect -125 -4878 -33 -4872
rect 33 -4838 125 -4832
rect 33 -4872 45 -4838
rect 113 -4872 125 -4838
rect 33 -4878 125 -4872
rect 191 -4838 283 -4832
rect 191 -4872 203 -4838
rect 271 -4872 283 -4838
rect 191 -4878 283 -4872
rect 349 -4838 441 -4832
rect 349 -4872 361 -4838
rect 429 -4872 441 -4838
rect 349 -4878 441 -4872
<< properties >>
string gencell sky130_fd_pr__nfet_03v3_nvt
string FIXED_BBOX -608 -4993 608 4993
string parameters w 48 l 0.50 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
