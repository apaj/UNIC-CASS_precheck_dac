magic
tech sky130A
magscale 1 2
timestamp 1695142129
<< dnwell >>
rect -1168 -5937 1168 5937
<< nwell >>
rect -1248 5731 1248 6017
rect -1248 -5731 -962 5731
rect 962 -5731 1248 5731
rect -1248 -6017 1248 -5731
<< pwell >>
rect -962 5573 -140 5731
rect -962 115 -140 273
rect 140 5573 962 5731
rect 140 115 962 273
rect -962 -273 -140 -115
rect -962 -5731 -140 -5573
rect 140 -273 962 -115
rect 140 -5731 962 -5573
<< rpw >>
rect -962 273 -140 5573
rect 140 273 962 5573
rect -962 -5573 -140 -273
rect 140 -5573 962 -273
<< psubdiff >>
rect -922 5573 -898 5679
rect -204 5573 -180 5679
rect 180 5573 204 5679
rect 898 5573 922 5679
rect -922 167 -898 273
rect -204 167 -180 273
rect 180 167 204 273
rect 898 167 922 273
rect -922 -273 -898 -167
rect -204 -273 -180 -167
rect 180 -273 204 -167
rect 898 -273 922 -167
rect -922 -5679 -898 -5573
rect -204 -5679 -180 -5573
rect 180 -5679 204 -5573
rect 898 -5679 922 -5573
<< nsubdiff >>
rect -1122 5857 -1026 5891
rect 1026 5857 1122 5891
rect -1122 5795 -1088 5857
rect 1088 5795 1122 5857
rect -1122 -5857 -1088 -5795
rect 1088 -5857 1122 -5795
rect -1122 -5891 -1026 -5857
rect 1026 -5891 1122 -5857
<< psubdiffcont >>
rect -898 5573 -204 5679
rect 204 5573 898 5679
rect -898 167 -204 273
rect 204 167 898 273
rect -898 -273 -204 -167
rect 204 -273 898 -167
rect -898 -5679 -204 -5573
rect 204 -5679 898 -5573
<< nsubdiffcont >>
rect -1026 5857 1026 5891
rect -1122 -5795 -1088 5795
rect 1088 -5795 1122 5795
rect -1026 -5891 1026 -5857
<< locali >>
rect -1122 5857 -1026 5891
rect 1026 5857 1122 5891
rect -1122 5795 -1088 5857
rect 1088 5795 1122 5857
rect -914 5643 -898 5679
rect -204 5643 -188 5679
rect -914 5590 -910 5643
rect -192 5590 -188 5643
rect -914 5573 -898 5590
rect -204 5573 -188 5590
rect 188 5643 204 5679
rect 898 5643 914 5679
rect 188 5590 192 5643
rect 910 5590 914 5643
rect 188 5573 204 5590
rect 898 5573 914 5590
rect -914 256 -898 273
rect -204 256 -188 273
rect -914 203 -910 256
rect -192 203 -188 256
rect -914 167 -898 203
rect -204 167 -188 203
rect 188 256 204 273
rect 898 256 914 273
rect 188 203 192 256
rect 910 203 914 256
rect 188 167 204 203
rect 898 167 914 203
rect -914 -203 -898 -167
rect -204 -203 -188 -167
rect -914 -256 -910 -203
rect -192 -256 -188 -203
rect -914 -273 -898 -256
rect -204 -273 -188 -256
rect 188 -203 204 -167
rect 898 -203 914 -167
rect 188 -256 192 -203
rect 910 -256 914 -203
rect 188 -273 204 -256
rect 898 -273 914 -256
rect -914 -5590 -898 -5573
rect -204 -5590 -188 -5573
rect -914 -5643 -910 -5590
rect -192 -5643 -188 -5590
rect -914 -5679 -898 -5643
rect -204 -5679 -188 -5643
rect 188 -5590 204 -5573
rect 898 -5590 914 -5573
rect 188 -5643 192 -5590
rect 910 -5643 914 -5590
rect 188 -5679 204 -5643
rect 898 -5679 914 -5643
rect -1122 -5857 -1088 -5795
rect 1088 -5857 1122 -5795
rect -1122 -5891 -1026 -5857
rect 1026 -5891 1122 -5857
<< viali >>
rect -910 5590 -898 5643
rect -898 5590 -204 5643
rect -204 5590 -192 5643
rect 192 5590 204 5643
rect 204 5590 898 5643
rect 898 5590 910 5643
rect -910 203 -898 256
rect -898 203 -204 256
rect -204 203 -192 256
rect 192 203 204 256
rect 204 203 898 256
rect 898 203 910 256
rect -910 -256 -898 -203
rect -898 -256 -204 -203
rect -204 -256 -192 -203
rect 192 -256 204 -203
rect 204 -256 898 -203
rect 898 -256 910 -203
rect -910 -5643 -898 -5590
rect -898 -5643 -204 -5590
rect -204 -5643 -192 -5590
rect 192 -5643 204 -5590
rect 204 -5643 898 -5590
rect 898 -5643 910 -5590
<< metal1 >>
rect -922 5643 -180 5649
rect -922 5590 -910 5643
rect -192 5590 -180 5643
rect -922 5584 -180 5590
rect 180 5643 922 5649
rect 180 5590 192 5643
rect 910 5590 922 5643
rect 180 5584 922 5590
rect -922 256 -180 262
rect -922 203 -910 256
rect -192 203 -180 256
rect -922 197 -180 203
rect 180 256 922 262
rect 180 203 192 256
rect 910 203 922 256
rect 180 197 922 203
rect -922 -203 -180 -197
rect -922 -256 -910 -203
rect -192 -256 -180 -203
rect -922 -262 -180 -256
rect 180 -203 922 -197
rect 180 -256 192 -203
rect 910 -256 922 -203
rect 180 -262 922 -256
rect -922 -5590 -180 -5584
rect -922 -5643 -910 -5590
rect -192 -5643 -180 -5590
rect -922 -5649 -180 -5643
rect 180 -5590 922 -5584
rect 180 -5643 192 -5590
rect 910 -5643 922 -5590
rect 180 -5649 922 -5643
<< properties >>
string FIXED_BBOX -1105 -5874 1105 5874
string gencell sky130_fd_pr__res_iso_pw
string library sky130
string parameters w 4.110 l 26.50 m 2 nx 2 wmin 2.650 lmin 26.50 rho 975 val 6.694k dummy 0 dw 0.25 term 1.0 guard 1 endcov 100 full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
