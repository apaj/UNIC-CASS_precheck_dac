magic
tech sky130A
magscale 1 2
timestamp 1697704145
<< nwell >>
rect 2166 2774 2472 3562
rect 2448 1014 3188 1368
<< viali >>
rect 3790 5544 3830 5750
rect 3788 5056 3828 5262
rect 3794 4584 3834 4790
rect 984 4388 1156 4536
rect 3788 4104 3828 4310
rect 1624 2854 1996 2894
rect 2288 2334 2484 2570
rect 3506 2314 3764 2580
rect 2644 1446 3016 1486
rect 2618 902 2990 942
rect 3898 910 4220 946
rect 2198 -232 2456 20
<< metal1 >>
rect 3764 5762 3846 5770
rect 3764 5750 3970 5762
rect -278 5538 -78 5540
rect 1564 5538 1990 5714
rect -278 5340 1990 5538
rect 146 5314 1990 5340
rect 146 3260 438 5314
rect 1564 5100 1990 5314
rect 1570 4570 1996 4762
rect 920 4536 1996 4570
rect 920 4388 984 4536
rect 1156 4388 1996 4536
rect 920 4356 1996 4388
rect 1570 4148 1996 4356
rect 3264 4148 3712 5714
rect 3764 5544 3790 5750
rect 3830 5544 3970 5750
rect 3764 5262 3970 5544
rect 3764 5056 3788 5262
rect 3828 5056 3970 5262
rect 3764 4790 3970 5056
rect 3764 4584 3794 4790
rect 3834 4584 3970 4790
rect 3764 4310 3970 4584
rect 3764 4120 3788 4310
rect 3762 4104 3788 4120
rect 3828 4104 3970 4310
rect 3762 3866 3970 4104
rect 1722 3592 2920 3720
rect 3762 3674 3962 3866
rect 1724 3322 1896 3592
rect 2240 3274 2424 3592
rect 2744 3316 2916 3592
rect 146 3082 1698 3260
rect 1920 3218 2424 3274
rect 1920 3084 2428 3218
rect 146 2944 398 3082
rect 2232 2958 2428 3084
rect 146 2894 2016 2944
rect 146 2854 1624 2894
rect 1996 2854 2016 2894
rect 146 2842 2016 2854
rect 1592 1532 2016 2842
rect 2232 2762 2436 2958
rect 2236 2758 2436 2762
rect 2202 2570 2696 2648
rect 2202 2334 2288 2570
rect 2484 2334 2696 2570
rect 2202 2240 2696 2334
rect 2944 2580 3834 2660
rect 2944 2314 3506 2580
rect 3764 2314 3834 2580
rect 2944 2248 3834 2314
rect 1588 1486 3038 1532
rect 1588 1446 2644 1486
rect 3016 1446 3038 1486
rect 1588 1418 3038 1446
rect 2610 982 3018 1418
rect 2610 946 4230 982
rect 2610 942 3898 946
rect 2610 902 2618 942
rect 2990 910 3898 942
rect 4220 910 4230 946
rect 2990 902 4230 910
rect 2610 876 4230 902
rect 2612 874 4230 876
rect 2150 20 2684 194
rect 3100 158 3320 162
rect 2150 -232 2198 20
rect 2456 -232 2684 20
rect 2150 -392 2684 -232
rect 2920 -342 3320 158
rect 3366 28 3936 190
rect 4326 178 4574 182
rect 3366 -222 3394 28
rect 3604 -222 3936 28
rect 3366 -300 3936 -222
rect 4146 -322 4574 178
rect 2712 -1546 2896 -922
rect 3100 -1406 3320 -342
rect 3130 -1482 3320 -1406
rect 2708 -1732 2898 -1546
rect 3126 -1682 3326 -1482
rect 3948 -1576 4132 -906
rect 4326 -1386 4574 -322
rect 3944 -1642 4132 -1576
rect 4378 -1448 4574 -1386
rect 2706 -1932 2906 -1732
rect 3944 -1842 4146 -1642
rect 4378 -1648 4578 -1448
<< via1 >>
rect 984 4388 1156 4536
rect 2288 2334 2484 2570
rect 3506 2314 3764 2580
rect 2198 -232 2456 20
rect 3394 -222 3604 28
<< metal2 >>
rect 882 4536 1238 4572
rect 882 4388 984 4536
rect 1156 4388 1238 4536
rect 882 2616 1238 4388
rect 882 2570 2602 2616
rect 882 2334 2288 2570
rect 2484 2334 2602 2570
rect 882 2278 2602 2334
rect 1012 2274 2602 2278
rect 3450 2580 3862 2660
rect 3450 2314 3506 2580
rect 3764 2360 3862 2580
rect 3764 2314 3866 2360
rect 3450 1288 3866 2314
rect 2150 1130 3866 1288
rect 2150 1128 3616 1130
rect 2154 94 2484 1128
rect 2142 20 2500 94
rect 2142 -232 2198 20
rect 2456 -232 2500 20
rect 2142 -298 2500 -232
rect 3366 28 3616 1128
rect 3366 -222 3394 28
rect 3604 -222 3616 28
rect 3366 -274 3616 -222
use sky130_fd_pr__pfet_g5v0d10v5_FGUWVM  XM1
timestamp 1697704145
transform 1 0 1808 0 1 3171
box -358 -397 358 397
use sky130_fd_pr__pfet_g5v0d10v5_FG5HVM  XM2
timestamp 1697704145
transform 1 0 2830 0 1 2465
box -358 -1097 358 1097
use sky130_fd_pr__pfet_g5v0d10v5_FG5HVM  XM3
timestamp 1697704145
transform 1 0 2806 0 1 -83
box -358 -1097 358 1097
use sky130_fd_pr__pfet_g5v0d10v5_FG5HVM  XM4
timestamp 1697704145
transform 1 0 4038 0 1 -79
box -358 -1097 358 1097
use sky130_fd_pr__res_xhigh_po_0p69_C4MSH5  XR1
timestamp 1697704145
transform 0 -1 2636 1 0 4207
box -235 -1228 235 1228
use sky130_fd_pr__res_xhigh_po_0p69_C4MSH5  XR2
timestamp 1697704145
transform 0 -1 2636 1 0 4687
box -235 -1228 235 1228
use sky130_fd_pr__res_xhigh_po_0p69_C4MSH5  XR3
timestamp 1697704145
transform 0 -1 2636 1 0 5161
box -235 -1228 235 1228
use sky130_fd_pr__res_xhigh_po_0p69_C4MSH5  XR4
timestamp 1697704145
transform 0 -1 2634 1 0 5643
box -235 -1228 235 1228
<< labels >>
flabel metal1 -278 5340 -78 5540 0 FreeSans 1280 0 0 0 vsup
port 0 nsew
flabel metal1 3762 3674 3962 3874 0 FreeSans 1280 0 0 0 vgnd
port 1 nsew
flabel metal1 2236 2758 2436 2958 0 FreeSans 1280 0 0 0 iref
port 2 nsew
flabel metal1 3126 -1682 3326 -1482 0 FreeSans 1280 0 0 0 iout
port 4 nsew
flabel metal1 2706 -1932 2906 -1732 0 FreeSans 1280 0 0 0 vsw
port 3 nsew
flabel metal1 3946 -1842 4146 -1642 0 FreeSans 1280 0 0 0 vbias
port 6 nsew
flabel metal1 4378 -1648 4578 -1448 0 FreeSans 1280 0 0 0 iout_n
port 5 nsew
rlabel metal1 3348 4624 3560 5140 1 parR
rlabel metal2 3586 1336 3798 1852 1 sourceM3M4
rlabel metal2 936 3524 1148 4040 1 sourceM2
<< end >>
