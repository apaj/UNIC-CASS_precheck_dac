magic
tech sky130A
magscale 1 2
timestamp 1697619488
<< viali >>
rect -1516 4324 -1438 4396
<< metal1 >>
rect -1922 9024 -1718 10290
rect 1374 9100 6792 9172
rect -1922 8882 -834 9024
rect -1306 8632 -1232 8790
rect -1838 8400 -844 8538
rect -1826 7974 -1674 8400
rect 360 8394 782 9030
rect 1332 8976 6680 8982
rect 1332 8716 1350 8976
rect 1402 8974 6680 8976
rect 1402 8716 1620 8974
rect 1332 8714 1620 8716
rect 1672 8714 1900 8974
rect 1952 8714 2174 8974
rect 2226 8714 2454 8974
rect 2506 8714 2732 8974
rect 2784 8714 3010 8974
rect 3062 8714 3290 8974
rect 3342 8714 3566 8974
rect 3618 8714 3844 8974
rect 3896 8714 4122 8974
rect 4174 8714 4400 8974
rect 4452 8714 4678 8974
rect 4730 8714 4956 8974
rect 5008 8714 5234 8974
rect 5286 8714 5512 8974
rect 5564 8714 5788 8974
rect 5840 8714 6068 8974
rect 6120 8714 6346 8974
rect 6398 8714 6622 8974
rect 6674 8714 6680 8974
rect 1332 8706 6680 8714
rect 1458 8498 6842 8504
rect 1458 8492 2056 8498
rect 1458 8478 1774 8492
rect -1590 8268 -1070 8304
rect 1458 8218 1502 8478
rect 1554 8232 1774 8478
rect 1826 8238 2056 8492
rect 2108 8496 6842 8498
rect 2108 8238 2332 8496
rect 1826 8236 2332 8238
rect 2384 8236 2610 8496
rect 2662 8236 2890 8496
rect 2942 8236 3166 8496
rect 3218 8236 3446 8496
rect 3498 8236 3722 8496
rect 3774 8236 4000 8496
rect 4052 8236 4278 8496
rect 4330 8236 4556 8496
rect 4608 8236 4836 8496
rect 4888 8236 5112 8496
rect 5164 8236 5392 8496
rect 5444 8236 5668 8496
rect 5720 8236 5946 8496
rect 5998 8236 6226 8496
rect 6278 8236 6502 8496
rect 6554 8236 6780 8496
rect 6832 8236 6842 8496
rect 1826 8232 6842 8236
rect 1554 8218 6842 8232
rect 1458 8208 6842 8218
rect -1208 7916 -550 7956
rect -34 7912 622 7952
rect -1264 7770 -646 7776
rect -1264 7508 -1258 7770
rect -1206 7508 -982 7770
rect -930 7508 -704 7770
rect -652 7508 -646 7770
rect -1264 7502 -646 7508
rect -90 7770 526 7776
rect -90 7750 190 7770
rect -90 7490 -88 7750
rect -36 7510 190 7750
rect 242 7510 468 7770
rect 520 7510 526 7770
rect -36 7490 526 7510
rect -90 7484 526 7490
rect -1104 6934 -488 6940
rect -1104 6932 -546 6934
rect -1104 6670 -1098 6932
rect -1046 6670 -824 6932
rect -772 6672 -546 6932
rect -494 6672 -488 6934
rect -772 6670 -488 6672
rect -1104 6664 -488 6670
rect 62 6916 684 6922
rect 62 6656 68 6916
rect 120 6656 346 6916
rect 398 6656 626 6916
rect 678 6656 684 6916
rect 62 6650 684 6656
rect -1586 6080 -1552 6420
rect -1222 6382 -530 6432
rect -54 6380 638 6430
rect 1392 6382 6782 6432
rect -1314 6244 2302 6298
rect -1674 6018 2754 6080
rect -1342 5978 -1256 5984
rect -1342 5948 -1336 5978
rect -1494 5922 -1336 5948
rect -1264 5948 -1256 5978
rect -1264 5922 -1090 5948
rect -1494 5900 -1090 5922
rect 526 5878 2586 5926
rect -694 5828 -624 5834
rect -1544 5814 -1198 5820
rect -1544 5554 -1538 5814
rect -1482 5554 -1260 5814
rect -1204 5554 -1198 5814
rect -694 5568 -688 5828
rect -630 5568 -624 5828
rect -694 5562 -624 5568
rect -128 5820 -58 5826
rect -128 5560 -122 5820
rect -64 5560 -58 5820
rect -128 5554 -58 5560
rect 462 5806 2486 5816
rect -1544 5548 -1198 5554
rect 462 5546 474 5806
rect 530 5546 752 5806
rect 808 5546 1028 5806
rect 1084 5546 1306 5806
rect 1362 5546 1584 5806
rect 1640 5546 1864 5806
rect 1920 5546 2142 5806
rect 2198 5546 2420 5806
rect 2476 5546 2486 5806
rect 462 5538 2486 5546
rect -536 5234 -466 5240
rect -1386 5224 -1040 5230
rect -1386 4964 -1380 5224
rect -1324 4964 -1102 5224
rect -1046 4964 -1040 5224
rect -536 4972 -530 5234
rect -472 4972 -466 5234
rect -536 4966 -466 4972
rect 30 5234 100 5240
rect 30 4972 36 5234
rect 94 4972 100 5234
rect 30 4966 100 4972
rect 624 5014 2640 5020
rect -1386 4958 -1040 4964
rect -3490 4738 -2778 4856
rect -1484 4788 -1106 4836
rect -624 4828 -540 4830
rect -3490 4444 -3170 4738
rect -2876 4444 -2778 4738
rect -3490 4438 -2778 4444
rect -3488 4436 -3288 4438
rect -1328 4414 -1252 4788
rect -624 4762 -614 4828
rect -544 4762 -540 4828
rect -624 4734 -540 4762
rect -466 4822 -378 4824
rect -466 4778 36 4822
rect -1020 4700 -930 4704
rect -1020 4648 -1008 4700
rect -944 4698 -930 4700
rect -944 4696 -682 4698
rect -466 4696 -378 4778
rect 624 4754 630 5014
rect 688 4754 908 5014
rect 966 4754 1186 5014
rect 1244 4754 1464 5014
rect 1522 4754 1742 5014
rect 1800 4754 2020 5014
rect 2078 4754 2298 5014
rect 2356 4754 2576 5014
rect 2634 4754 2640 5014
rect 624 4748 2640 4754
rect -944 4672 -378 4696
rect -944 4648 -380 4672
rect -1020 4646 -380 4648
rect -1020 4640 -930 4646
rect -718 4644 -380 4646
rect -126 4512 -20 4678
rect 526 4568 2576 4614
rect -2218 4406 -2076 4410
rect -2218 4402 -1556 4406
rect -2218 4396 -1420 4402
rect -2218 4324 -1516 4396
rect -1438 4324 -1420 4396
rect -1328 4372 -100 4414
rect -2218 4312 -1420 4324
rect -2218 3984 -2076 4312
rect -542 4280 -196 4286
rect -542 4020 -536 4280
rect -480 4020 -258 4280
rect -202 4020 -196 4280
rect -542 4014 -196 4020
rect -3488 3980 -2076 3984
rect -3496 3782 -2076 3980
rect -3496 3780 -2190 3782
rect -382 3636 -38 3642
rect -382 3634 -100 3636
rect -382 3374 -376 3634
rect -320 3376 -100 3634
rect -44 3376 -38 3636
rect -320 3374 -38 3376
rect -382 3368 -38 3374
rect -1880 2630 -1628 2648
rect -1880 2468 -1850 2630
rect -1640 2468 -1628 2630
rect -1880 2212 -1628 2468
rect 0 -800 200 -600
<< via1 >>
rect 1350 8716 1402 8976
rect 1620 8714 1672 8974
rect 1900 8714 1952 8974
rect 2174 8714 2226 8974
rect 2454 8714 2506 8974
rect 2732 8714 2784 8974
rect 3010 8714 3062 8974
rect 3290 8714 3342 8974
rect 3566 8714 3618 8974
rect 3844 8714 3896 8974
rect 4122 8714 4174 8974
rect 4400 8714 4452 8974
rect 4678 8714 4730 8974
rect 4956 8714 5008 8974
rect 5234 8714 5286 8974
rect 5512 8714 5564 8974
rect 5788 8714 5840 8974
rect 6068 8714 6120 8974
rect 6346 8714 6398 8974
rect 6622 8714 6674 8974
rect 1502 8218 1554 8478
rect 1774 8232 1826 8492
rect 2056 8238 2108 8498
rect 2332 8236 2384 8496
rect 2610 8236 2662 8496
rect 2890 8236 2942 8496
rect 3166 8236 3218 8496
rect 3446 8236 3498 8496
rect 3722 8236 3774 8496
rect 4000 8236 4052 8496
rect 4278 8236 4330 8496
rect 4556 8236 4608 8496
rect 4836 8236 4888 8496
rect 5112 8236 5164 8496
rect 5392 8236 5444 8496
rect 5668 8236 5720 8496
rect 5946 8236 5998 8496
rect 6226 8236 6278 8496
rect 6502 8236 6554 8496
rect 6780 8236 6832 8496
rect -1258 7508 -1206 7770
rect -982 7508 -930 7770
rect -704 7508 -652 7770
rect -88 7490 -36 7750
rect 190 7510 242 7770
rect 468 7510 520 7770
rect -1804 6366 -1706 6682
rect -1098 6670 -1046 6932
rect -824 6670 -772 6932
rect -546 6672 -494 6934
rect 68 6656 120 6916
rect 346 6656 398 6916
rect 626 6656 678 6916
rect -1336 5922 -1264 5978
rect -1538 5554 -1482 5814
rect -1260 5554 -1204 5814
rect -688 5568 -630 5828
rect -122 5560 -64 5820
rect 474 5546 530 5806
rect 752 5546 808 5806
rect 1028 5546 1084 5806
rect 1306 5546 1362 5806
rect 1584 5546 1640 5806
rect 1864 5546 1920 5806
rect 2142 5546 2198 5806
rect 2420 5546 2476 5806
rect -1380 4964 -1324 5224
rect -1102 4964 -1046 5224
rect -530 4972 -472 5234
rect 36 4972 94 5234
rect -3170 4444 -2876 4738
rect -614 4762 -544 4828
rect -1008 4648 -944 4700
rect 630 4754 688 5014
rect 908 4754 966 5014
rect 1186 4754 1244 5014
rect 1464 4754 1522 5014
rect 1742 4754 1800 5014
rect 2020 4754 2078 5014
rect 2298 4754 2356 5014
rect 2576 4754 2634 5014
rect -536 4020 -480 4280
rect -258 4020 -202 4280
rect -376 3374 -320 3634
rect -100 3376 -44 3636
rect -1850 2468 -1640 2630
<< metal2 >>
rect 1332 8976 6680 8982
rect 1332 8716 1350 8976
rect 1402 8974 6680 8976
rect 1402 8716 1620 8974
rect 1332 8714 1620 8716
rect 1672 8714 1900 8974
rect 1952 8714 2174 8974
rect 2226 8714 2454 8974
rect 2506 8714 2732 8974
rect 2784 8714 3010 8974
rect 3062 8714 3290 8974
rect 3342 8714 3566 8974
rect 3618 8714 3844 8974
rect 3896 8714 4122 8974
rect 4174 8714 4400 8974
rect 4452 8714 4678 8974
rect 4730 8714 4956 8974
rect 5008 8714 5234 8974
rect 5286 8714 5512 8974
rect 5564 8714 5788 8974
rect 5840 8714 6068 8974
rect 6120 8714 6346 8974
rect 6398 8714 6622 8974
rect 6674 8714 6680 8974
rect 1332 8706 6680 8714
rect 1458 8498 6842 8504
rect 1458 8492 2056 8498
rect 1458 8478 1774 8492
rect 1458 8218 1502 8478
rect 1554 8232 1774 8478
rect 1826 8238 2056 8492
rect 2108 8496 6842 8498
rect 2108 8238 2332 8496
rect 1826 8236 2332 8238
rect 2384 8236 2610 8496
rect 2662 8236 2890 8496
rect 2942 8236 3166 8496
rect 3218 8236 3446 8496
rect 3498 8236 3722 8496
rect 3774 8236 4000 8496
rect 4052 8236 4278 8496
rect 4330 8236 4556 8496
rect 4608 8236 4836 8496
rect 4888 8236 5112 8496
rect 5164 8236 5392 8496
rect 5444 8236 5668 8496
rect 5720 8236 5946 8496
rect 5998 8236 6226 8496
rect 6278 8236 6502 8496
rect 6554 8236 6780 8496
rect 6832 8236 6842 8496
rect 1826 8232 6842 8236
rect 1554 8218 6842 8232
rect 1458 8208 6842 8218
rect -1264 7770 -646 7776
rect -1264 7508 -1258 7770
rect -1206 7508 -982 7770
rect -930 7508 -704 7770
rect -652 7508 -646 7770
rect -1264 7502 -646 7508
rect -90 7770 526 7776
rect -90 7750 190 7770
rect -90 7490 -88 7750
rect -36 7510 190 7750
rect 242 7510 468 7770
rect 520 7510 526 7770
rect -36 7490 526 7510
rect -90 7484 526 7490
rect -1104 6934 -488 6940
rect -1104 6932 -546 6934
rect -1852 6682 -1658 6736
rect -1852 6366 -1804 6682
rect -1706 6366 -1658 6682
rect -1104 6670 -1098 6932
rect -1046 6670 -824 6932
rect -772 6672 -546 6932
rect -494 6672 -488 6934
rect -772 6670 -488 6672
rect -1104 6664 -488 6670
rect 62 6916 684 6922
rect 62 6656 68 6916
rect 120 6656 346 6916
rect 398 6656 626 6916
rect 678 6656 684 6916
rect 62 6650 684 6656
rect -1852 6348 -1658 6366
rect -1852 6118 -1656 6348
rect -1102 6146 -1048 6148
rect -1328 6118 -1048 6146
rect -1852 6038 -1252 6118
rect -1816 6036 -1252 6038
rect -1346 5978 -1254 6036
rect -1346 5922 -1336 5978
rect -1264 5922 -1254 5978
rect -1346 5916 -1254 5922
rect -1544 5814 -1198 5820
rect -1544 5764 -1538 5814
rect -1974 5570 -1538 5764
rect -3230 4742 -2682 4924
rect -3230 4738 -3146 4742
rect -3230 4444 -3170 4738
rect -3230 4380 -3146 4444
rect -2790 4380 -2682 4742
rect -3230 4188 -2682 4380
rect -1974 4282 -1764 5570
rect -1544 5554 -1538 5570
rect -1482 5554 -1260 5814
rect -1204 5554 -1198 5814
rect -1544 5548 -1198 5554
rect -1102 5230 -1048 6118
rect -694 5828 -624 5834
rect -694 5568 -688 5828
rect -630 5826 -64 5828
rect -630 5820 -58 5826
rect -630 5572 -122 5820
rect -630 5568 -624 5572
rect -694 5562 -624 5568
rect -536 5234 -466 5240
rect -1386 5224 -1040 5230
rect -1386 4964 -1380 5224
rect -1324 4964 -1102 5224
rect -1046 4964 -1040 5224
rect -536 4972 -530 5234
rect -472 4972 -466 5234
rect -536 4966 -466 4972
rect -1386 4958 -1040 4964
rect -624 4828 -534 4838
rect -624 4762 -614 4828
rect -544 4762 -534 4828
rect -1482 4700 -930 4712
rect -1482 4648 -1008 4700
rect -944 4648 -930 4700
rect -1482 4640 -930 4648
rect -1482 4422 -1400 4640
rect -624 4558 -534 4762
rect -364 4648 -228 5572
rect -128 5560 -122 5572
rect -64 5560 -58 5820
rect -128 5554 -58 5560
rect 462 5806 2486 5816
rect 462 5546 474 5806
rect 530 5546 752 5806
rect 808 5546 1028 5806
rect 1084 5546 1306 5806
rect 1362 5546 1584 5806
rect 1640 5546 1864 5806
rect 1920 5546 2142 5806
rect 2198 5546 2420 5806
rect 2476 5546 2486 5806
rect 462 5538 2486 5546
rect 30 5234 100 5240
rect 30 4972 36 5234
rect 94 4972 100 5234
rect 30 4966 100 4972
rect 624 5014 2640 5020
rect 624 4754 630 5014
rect 688 4754 908 5014
rect 966 4754 1186 5014
rect 1244 4754 1464 5014
rect 1522 4754 1742 5014
rect 1800 4754 2020 5014
rect 2078 4754 2298 5014
rect 2356 4754 2576 5014
rect 2634 4754 2640 5014
rect 624 4748 2640 4754
rect -364 4568 214 4648
rect -344 4558 214 4568
rect -920 4546 -534 4558
rect -920 4466 -908 4546
rect -806 4466 -534 4546
rect -920 4454 -534 4466
rect -1522 4320 -1398 4422
rect -542 4282 -196 4286
rect -1974 4280 -196 4282
rect -1974 4022 -536 4280
rect -1974 2686 -1764 4022
rect -542 4020 -536 4022
rect -480 4020 -258 4280
rect -202 4020 -196 4280
rect -542 4014 -196 4020
rect -382 3636 -38 3642
rect 78 3636 208 4558
rect -382 3634 -100 3636
rect -382 3374 -376 3634
rect -320 3376 -100 3634
rect -44 3388 210 3636
rect -44 3376 -38 3388
rect -320 3374 -38 3376
rect -382 3368 -38 3374
rect -1974 2630 -1564 2686
rect -1974 2468 -1850 2630
rect -1640 2468 -1564 2630
rect -1974 2462 -1564 2468
rect -1884 2454 -1564 2462
<< via2 >>
rect -3146 4738 -2790 4742
rect -3146 4444 -2876 4738
rect -2876 4444 -2790 4738
rect -3146 4380 -2790 4444
rect -908 4466 -806 4546
<< metal3 >>
rect -3176 4742 -2772 4774
rect -3176 4380 -3146 4742
rect -2790 4560 -2772 4742
rect -2790 4546 -794 4560
rect -2790 4466 -908 4546
rect -806 4466 -794 4546
rect -2790 4454 -794 4466
rect -2790 4380 -2772 4454
rect -3176 4360 -2772 4380
use sky130_fd_pr__cap_mim_m3_1_C5B489  XC1
timestamp 1697533315
transform 1 0 3962 0 1 4642
box -1150 -1500 1149 1500
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM1
timestamp 1697533315
transform 1 0 -580 0 1 5364
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM2
timestamp 1697533315
transform 1 0 -14 0 1 5356
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_NQCFE9  XM3
timestamp 1697536037
transform 1 0 -1293 0 1 5364
box -417 -758 417 758
use sky130_fd_pr__nfet_g5v0d10v5_CJGAEC  XM4
timestamp 1697536037
transform 1 0 -289 0 1 3836
box -417 -758 417 758
use sky130_fd_pr__nfet_g5v0d10v5_2MGL8M  XM5
timestamp 1697536037
transform 1 0 1553 0 1 5246
box -1251 -858 1251 858
use sky130_fd_pr__pfet_g5v0d10v5_X3UTN5  XM6
timestamp 1697536037
transform 1 0 -876 0 1 7171
box -586 -997 586 997
use sky130_fd_pr__pfet_g5v0d10v5_AE43MT  XM7
timestamp 1697536280
transform 1 0 294 0 1 7169
box -586 -997 586 997
use sky130_fd_pr__pfet_g5v0d10v5_CNRWF7  XM8
timestamp 1697534501
transform 1 0 4087 0 1 7771
box -2949 -1597 2949 1597
use sky130_fd_pr__res_xhigh_po_0p69_5CVACY  XR1
timestamp 1697533315
transform 1 0 -1751 0 1 7372
box -235 -1198 235 1198
use sky130_fd_pr__res_xhigh_po_0p69_5CVACY  XR2
timestamp 1697533315
transform 0 -1 -240 1 0 8467
box -235 -1198 235 1198
use sky130_fd_pr__res_xhigh_po_0p69_5CVACY  XR3
timestamp 1697533315
transform 0 1 -244 -1 0 8955
box -235 -1198 235 1198
<< labels >>
flabel metal1 0 -800 200 -600 0 FreeSans 1280 0 0 0 outSingle
port 2 nsew
flabel metal1 -1920 10086 -1720 10286 0 FreeSans 1280 0 0 0 power
port 3 nsew
flabel metal1 -1880 2212 -1680 2412 0 FreeSans 1280 0 0 0 ground
port 4 nsew
flabel metal1 -3488 4436 -3288 4636 0 FreeSans 1280 0 0 0 inPos
port 0 nsew
flabel metal1 -3496 3780 -3296 3980 0 FreeSans 1280 0 0 0 inNeg
port 1 nsew
<< end >>
