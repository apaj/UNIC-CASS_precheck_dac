**.subckt dac_cell1 vsup vgnd iref vsw iout iout_n vbias
*.iopin vsup
*.iopin vgnd
*.iopin iref
*.iopin vsw
*.iopin iout
*.iopin iout_n
*.iopin vbias
XM1 iref iref vsup vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 sourceM3M4 iref sourceM2 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 iout vsw sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 iout_n vbias sourceM3M4 vsup sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XR1 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
XR2 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
XR3 parR vsup vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
XR4 sourceM2 parR vgnd sky130_fd_pr__res_xhigh_po_0p69 L=58 mult=1 m=1
**.ends
** flattened .save nodes
.end
