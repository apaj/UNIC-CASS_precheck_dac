magic
tech sky130A
magscale 1 2
timestamp 1697933062
<< nwell >>
rect -2949 -1597 2949 1597
<< mvpmos >>
rect -2691 -1300 -2591 1300
rect -2413 -1300 -2313 1300
rect -2135 -1300 -2035 1300
rect -1857 -1300 -1757 1300
rect -1579 -1300 -1479 1300
rect -1301 -1300 -1201 1300
rect -1023 -1300 -923 1300
rect -745 -1300 -645 1300
rect -467 -1300 -367 1300
rect -189 -1300 -89 1300
rect 89 -1300 189 1300
rect 367 -1300 467 1300
rect 645 -1300 745 1300
rect 923 -1300 1023 1300
rect 1201 -1300 1301 1300
rect 1479 -1300 1579 1300
rect 1757 -1300 1857 1300
rect 2035 -1300 2135 1300
rect 2313 -1300 2413 1300
rect 2591 -1300 2691 1300
<< mvpdiff >>
rect -2749 1288 -2691 1300
rect -2749 -1288 -2737 1288
rect -2703 -1288 -2691 1288
rect -2749 -1300 -2691 -1288
rect -2591 1288 -2533 1300
rect -2591 -1288 -2579 1288
rect -2545 -1288 -2533 1288
rect -2591 -1300 -2533 -1288
rect -2471 1288 -2413 1300
rect -2471 -1288 -2459 1288
rect -2425 -1288 -2413 1288
rect -2471 -1300 -2413 -1288
rect -2313 1288 -2255 1300
rect -2313 -1288 -2301 1288
rect -2267 -1288 -2255 1288
rect -2313 -1300 -2255 -1288
rect -2193 1288 -2135 1300
rect -2193 -1288 -2181 1288
rect -2147 -1288 -2135 1288
rect -2193 -1300 -2135 -1288
rect -2035 1288 -1977 1300
rect -2035 -1288 -2023 1288
rect -1989 -1288 -1977 1288
rect -2035 -1300 -1977 -1288
rect -1915 1288 -1857 1300
rect -1915 -1288 -1903 1288
rect -1869 -1288 -1857 1288
rect -1915 -1300 -1857 -1288
rect -1757 1288 -1699 1300
rect -1757 -1288 -1745 1288
rect -1711 -1288 -1699 1288
rect -1757 -1300 -1699 -1288
rect -1637 1288 -1579 1300
rect -1637 -1288 -1625 1288
rect -1591 -1288 -1579 1288
rect -1637 -1300 -1579 -1288
rect -1479 1288 -1421 1300
rect -1479 -1288 -1467 1288
rect -1433 -1288 -1421 1288
rect -1479 -1300 -1421 -1288
rect -1359 1288 -1301 1300
rect -1359 -1288 -1347 1288
rect -1313 -1288 -1301 1288
rect -1359 -1300 -1301 -1288
rect -1201 1288 -1143 1300
rect -1201 -1288 -1189 1288
rect -1155 -1288 -1143 1288
rect -1201 -1300 -1143 -1288
rect -1081 1288 -1023 1300
rect -1081 -1288 -1069 1288
rect -1035 -1288 -1023 1288
rect -1081 -1300 -1023 -1288
rect -923 1288 -865 1300
rect -923 -1288 -911 1288
rect -877 -1288 -865 1288
rect -923 -1300 -865 -1288
rect -803 1288 -745 1300
rect -803 -1288 -791 1288
rect -757 -1288 -745 1288
rect -803 -1300 -745 -1288
rect -645 1288 -587 1300
rect -645 -1288 -633 1288
rect -599 -1288 -587 1288
rect -645 -1300 -587 -1288
rect -525 1288 -467 1300
rect -525 -1288 -513 1288
rect -479 -1288 -467 1288
rect -525 -1300 -467 -1288
rect -367 1288 -309 1300
rect -367 -1288 -355 1288
rect -321 -1288 -309 1288
rect -367 -1300 -309 -1288
rect -247 1288 -189 1300
rect -247 -1288 -235 1288
rect -201 -1288 -189 1288
rect -247 -1300 -189 -1288
rect -89 1288 -31 1300
rect -89 -1288 -77 1288
rect -43 -1288 -31 1288
rect -89 -1300 -31 -1288
rect 31 1288 89 1300
rect 31 -1288 43 1288
rect 77 -1288 89 1288
rect 31 -1300 89 -1288
rect 189 1288 247 1300
rect 189 -1288 201 1288
rect 235 -1288 247 1288
rect 189 -1300 247 -1288
rect 309 1288 367 1300
rect 309 -1288 321 1288
rect 355 -1288 367 1288
rect 309 -1300 367 -1288
rect 467 1288 525 1300
rect 467 -1288 479 1288
rect 513 -1288 525 1288
rect 467 -1300 525 -1288
rect 587 1288 645 1300
rect 587 -1288 599 1288
rect 633 -1288 645 1288
rect 587 -1300 645 -1288
rect 745 1288 803 1300
rect 745 -1288 757 1288
rect 791 -1288 803 1288
rect 745 -1300 803 -1288
rect 865 1288 923 1300
rect 865 -1288 877 1288
rect 911 -1288 923 1288
rect 865 -1300 923 -1288
rect 1023 1288 1081 1300
rect 1023 -1288 1035 1288
rect 1069 -1288 1081 1288
rect 1023 -1300 1081 -1288
rect 1143 1288 1201 1300
rect 1143 -1288 1155 1288
rect 1189 -1288 1201 1288
rect 1143 -1300 1201 -1288
rect 1301 1288 1359 1300
rect 1301 -1288 1313 1288
rect 1347 -1288 1359 1288
rect 1301 -1300 1359 -1288
rect 1421 1288 1479 1300
rect 1421 -1288 1433 1288
rect 1467 -1288 1479 1288
rect 1421 -1300 1479 -1288
rect 1579 1288 1637 1300
rect 1579 -1288 1591 1288
rect 1625 -1288 1637 1288
rect 1579 -1300 1637 -1288
rect 1699 1288 1757 1300
rect 1699 -1288 1711 1288
rect 1745 -1288 1757 1288
rect 1699 -1300 1757 -1288
rect 1857 1288 1915 1300
rect 1857 -1288 1869 1288
rect 1903 -1288 1915 1288
rect 1857 -1300 1915 -1288
rect 1977 1288 2035 1300
rect 1977 -1288 1989 1288
rect 2023 -1288 2035 1288
rect 1977 -1300 2035 -1288
rect 2135 1288 2193 1300
rect 2135 -1288 2147 1288
rect 2181 -1288 2193 1288
rect 2135 -1300 2193 -1288
rect 2255 1288 2313 1300
rect 2255 -1288 2267 1288
rect 2301 -1288 2313 1288
rect 2255 -1300 2313 -1288
rect 2413 1288 2471 1300
rect 2413 -1288 2425 1288
rect 2459 -1288 2471 1288
rect 2413 -1300 2471 -1288
rect 2533 1288 2591 1300
rect 2533 -1288 2545 1288
rect 2579 -1288 2591 1288
rect 2533 -1300 2591 -1288
rect 2691 1288 2749 1300
rect 2691 -1288 2703 1288
rect 2737 -1288 2749 1288
rect 2691 -1300 2749 -1288
<< mvpdiffc >>
rect -2737 -1288 -2703 1288
rect -2579 -1288 -2545 1288
rect -2459 -1288 -2425 1288
rect -2301 -1288 -2267 1288
rect -2181 -1288 -2147 1288
rect -2023 -1288 -1989 1288
rect -1903 -1288 -1869 1288
rect -1745 -1288 -1711 1288
rect -1625 -1288 -1591 1288
rect -1467 -1288 -1433 1288
rect -1347 -1288 -1313 1288
rect -1189 -1288 -1155 1288
rect -1069 -1288 -1035 1288
rect -911 -1288 -877 1288
rect -791 -1288 -757 1288
rect -633 -1288 -599 1288
rect -513 -1288 -479 1288
rect -355 -1288 -321 1288
rect -235 -1288 -201 1288
rect -77 -1288 -43 1288
rect 43 -1288 77 1288
rect 201 -1288 235 1288
rect 321 -1288 355 1288
rect 479 -1288 513 1288
rect 599 -1288 633 1288
rect 757 -1288 791 1288
rect 877 -1288 911 1288
rect 1035 -1288 1069 1288
rect 1155 -1288 1189 1288
rect 1313 -1288 1347 1288
rect 1433 -1288 1467 1288
rect 1591 -1288 1625 1288
rect 1711 -1288 1745 1288
rect 1869 -1288 1903 1288
rect 1989 -1288 2023 1288
rect 2147 -1288 2181 1288
rect 2267 -1288 2301 1288
rect 2425 -1288 2459 1288
rect 2545 -1288 2579 1288
rect 2703 -1288 2737 1288
<< mvnsubdiff >>
rect -2883 1519 2883 1531
rect -2883 1485 -2775 1519
rect 2775 1485 2883 1519
rect -2883 1473 2883 1485
rect -2883 1423 -2825 1473
rect -2883 -1423 -2871 1423
rect -2837 -1423 -2825 1423
rect 2825 1423 2883 1473
rect -2883 -1473 -2825 -1423
rect 2825 -1423 2837 1423
rect 2871 -1423 2883 1423
rect 2825 -1473 2883 -1423
rect -2883 -1485 2883 -1473
rect -2883 -1519 -2775 -1485
rect 2775 -1519 2883 -1485
rect -2883 -1531 2883 -1519
<< mvnsubdiffcont >>
rect -2775 1485 2775 1519
rect -2871 -1423 -2837 1423
rect 2837 -1423 2871 1423
rect -2775 -1519 2775 -1485
<< poly >>
rect -2691 1381 -2591 1397
rect -2691 1347 -2675 1381
rect -2607 1347 -2591 1381
rect -2691 1300 -2591 1347
rect -2413 1381 -2313 1397
rect -2413 1347 -2397 1381
rect -2329 1347 -2313 1381
rect -2413 1300 -2313 1347
rect -2135 1381 -2035 1397
rect -2135 1347 -2119 1381
rect -2051 1347 -2035 1381
rect -2135 1300 -2035 1347
rect -1857 1381 -1757 1397
rect -1857 1347 -1841 1381
rect -1773 1347 -1757 1381
rect -1857 1300 -1757 1347
rect -1579 1381 -1479 1397
rect -1579 1347 -1563 1381
rect -1495 1347 -1479 1381
rect -1579 1300 -1479 1347
rect -1301 1381 -1201 1397
rect -1301 1347 -1285 1381
rect -1217 1347 -1201 1381
rect -1301 1300 -1201 1347
rect -1023 1381 -923 1397
rect -1023 1347 -1007 1381
rect -939 1347 -923 1381
rect -1023 1300 -923 1347
rect -745 1381 -645 1397
rect -745 1347 -729 1381
rect -661 1347 -645 1381
rect -745 1300 -645 1347
rect -467 1381 -367 1397
rect -467 1347 -451 1381
rect -383 1347 -367 1381
rect -467 1300 -367 1347
rect -189 1381 -89 1397
rect -189 1347 -173 1381
rect -105 1347 -89 1381
rect -189 1300 -89 1347
rect 89 1381 189 1397
rect 89 1347 105 1381
rect 173 1347 189 1381
rect 89 1300 189 1347
rect 367 1381 467 1397
rect 367 1347 383 1381
rect 451 1347 467 1381
rect 367 1300 467 1347
rect 645 1381 745 1397
rect 645 1347 661 1381
rect 729 1347 745 1381
rect 645 1300 745 1347
rect 923 1381 1023 1397
rect 923 1347 939 1381
rect 1007 1347 1023 1381
rect 923 1300 1023 1347
rect 1201 1381 1301 1397
rect 1201 1347 1217 1381
rect 1285 1347 1301 1381
rect 1201 1300 1301 1347
rect 1479 1381 1579 1397
rect 1479 1347 1495 1381
rect 1563 1347 1579 1381
rect 1479 1300 1579 1347
rect 1757 1381 1857 1397
rect 1757 1347 1773 1381
rect 1841 1347 1857 1381
rect 1757 1300 1857 1347
rect 2035 1381 2135 1397
rect 2035 1347 2051 1381
rect 2119 1347 2135 1381
rect 2035 1300 2135 1347
rect 2313 1381 2413 1397
rect 2313 1347 2329 1381
rect 2397 1347 2413 1381
rect 2313 1300 2413 1347
rect 2591 1381 2691 1397
rect 2591 1347 2607 1381
rect 2675 1347 2691 1381
rect 2591 1300 2691 1347
rect -2691 -1347 -2591 -1300
rect -2691 -1381 -2675 -1347
rect -2607 -1381 -2591 -1347
rect -2691 -1397 -2591 -1381
rect -2413 -1347 -2313 -1300
rect -2413 -1381 -2397 -1347
rect -2329 -1381 -2313 -1347
rect -2413 -1397 -2313 -1381
rect -2135 -1347 -2035 -1300
rect -2135 -1381 -2119 -1347
rect -2051 -1381 -2035 -1347
rect -2135 -1397 -2035 -1381
rect -1857 -1347 -1757 -1300
rect -1857 -1381 -1841 -1347
rect -1773 -1381 -1757 -1347
rect -1857 -1397 -1757 -1381
rect -1579 -1347 -1479 -1300
rect -1579 -1381 -1563 -1347
rect -1495 -1381 -1479 -1347
rect -1579 -1397 -1479 -1381
rect -1301 -1347 -1201 -1300
rect -1301 -1381 -1285 -1347
rect -1217 -1381 -1201 -1347
rect -1301 -1397 -1201 -1381
rect -1023 -1347 -923 -1300
rect -1023 -1381 -1007 -1347
rect -939 -1381 -923 -1347
rect -1023 -1397 -923 -1381
rect -745 -1347 -645 -1300
rect -745 -1381 -729 -1347
rect -661 -1381 -645 -1347
rect -745 -1397 -645 -1381
rect -467 -1347 -367 -1300
rect -467 -1381 -451 -1347
rect -383 -1381 -367 -1347
rect -467 -1397 -367 -1381
rect -189 -1347 -89 -1300
rect -189 -1381 -173 -1347
rect -105 -1381 -89 -1347
rect -189 -1397 -89 -1381
rect 89 -1347 189 -1300
rect 89 -1381 105 -1347
rect 173 -1381 189 -1347
rect 89 -1397 189 -1381
rect 367 -1347 467 -1300
rect 367 -1381 383 -1347
rect 451 -1381 467 -1347
rect 367 -1397 467 -1381
rect 645 -1347 745 -1300
rect 645 -1381 661 -1347
rect 729 -1381 745 -1347
rect 645 -1397 745 -1381
rect 923 -1347 1023 -1300
rect 923 -1381 939 -1347
rect 1007 -1381 1023 -1347
rect 923 -1397 1023 -1381
rect 1201 -1347 1301 -1300
rect 1201 -1381 1217 -1347
rect 1285 -1381 1301 -1347
rect 1201 -1397 1301 -1381
rect 1479 -1347 1579 -1300
rect 1479 -1381 1495 -1347
rect 1563 -1381 1579 -1347
rect 1479 -1397 1579 -1381
rect 1757 -1347 1857 -1300
rect 1757 -1381 1773 -1347
rect 1841 -1381 1857 -1347
rect 1757 -1397 1857 -1381
rect 2035 -1347 2135 -1300
rect 2035 -1381 2051 -1347
rect 2119 -1381 2135 -1347
rect 2035 -1397 2135 -1381
rect 2313 -1347 2413 -1300
rect 2313 -1381 2329 -1347
rect 2397 -1381 2413 -1347
rect 2313 -1397 2413 -1381
rect 2591 -1347 2691 -1300
rect 2591 -1381 2607 -1347
rect 2675 -1381 2691 -1347
rect 2591 -1397 2691 -1381
<< polycont >>
rect -2675 1347 -2607 1381
rect -2397 1347 -2329 1381
rect -2119 1347 -2051 1381
rect -1841 1347 -1773 1381
rect -1563 1347 -1495 1381
rect -1285 1347 -1217 1381
rect -1007 1347 -939 1381
rect -729 1347 -661 1381
rect -451 1347 -383 1381
rect -173 1347 -105 1381
rect 105 1347 173 1381
rect 383 1347 451 1381
rect 661 1347 729 1381
rect 939 1347 1007 1381
rect 1217 1347 1285 1381
rect 1495 1347 1563 1381
rect 1773 1347 1841 1381
rect 2051 1347 2119 1381
rect 2329 1347 2397 1381
rect 2607 1347 2675 1381
rect -2675 -1381 -2607 -1347
rect -2397 -1381 -2329 -1347
rect -2119 -1381 -2051 -1347
rect -1841 -1381 -1773 -1347
rect -1563 -1381 -1495 -1347
rect -1285 -1381 -1217 -1347
rect -1007 -1381 -939 -1347
rect -729 -1381 -661 -1347
rect -451 -1381 -383 -1347
rect -173 -1381 -105 -1347
rect 105 -1381 173 -1347
rect 383 -1381 451 -1347
rect 661 -1381 729 -1347
rect 939 -1381 1007 -1347
rect 1217 -1381 1285 -1347
rect 1495 -1381 1563 -1347
rect 1773 -1381 1841 -1347
rect 2051 -1381 2119 -1347
rect 2329 -1381 2397 -1347
rect 2607 -1381 2675 -1347
<< locali >>
rect -2871 1485 -2775 1519
rect 2775 1485 2871 1519
rect -2871 1423 -2837 1485
rect 2837 1423 2871 1485
rect -2691 1347 -2675 1381
rect -2607 1347 -2591 1381
rect -2413 1347 -2397 1381
rect -2329 1347 -2313 1381
rect -2135 1347 -2119 1381
rect -2051 1347 -2035 1381
rect -1857 1347 -1841 1381
rect -1773 1347 -1757 1381
rect -1579 1347 -1563 1381
rect -1495 1347 -1479 1381
rect -1301 1347 -1285 1381
rect -1217 1347 -1201 1381
rect -1023 1347 -1007 1381
rect -939 1347 -923 1381
rect -745 1347 -729 1381
rect -661 1347 -645 1381
rect -467 1347 -451 1381
rect -383 1347 -367 1381
rect -189 1347 -173 1381
rect -105 1347 -89 1381
rect 89 1347 105 1381
rect 173 1347 189 1381
rect 367 1347 383 1381
rect 451 1347 467 1381
rect 645 1347 661 1381
rect 729 1347 745 1381
rect 923 1347 939 1381
rect 1007 1347 1023 1381
rect 1201 1347 1217 1381
rect 1285 1347 1301 1381
rect 1479 1347 1495 1381
rect 1563 1347 1579 1381
rect 1757 1347 1773 1381
rect 1841 1347 1857 1381
rect 2035 1347 2051 1381
rect 2119 1347 2135 1381
rect 2313 1347 2329 1381
rect 2397 1347 2413 1381
rect 2591 1347 2607 1381
rect 2675 1347 2691 1381
rect -2737 1288 -2703 1304
rect -2737 -1304 -2703 -1288
rect -2579 1288 -2545 1304
rect -2579 -1304 -2545 -1288
rect -2459 1288 -2425 1304
rect -2459 -1304 -2425 -1288
rect -2301 1288 -2267 1304
rect -2301 -1304 -2267 -1288
rect -2181 1288 -2147 1304
rect -2181 -1304 -2147 -1288
rect -2023 1288 -1989 1304
rect -2023 -1304 -1989 -1288
rect -1903 1288 -1869 1304
rect -1903 -1304 -1869 -1288
rect -1745 1288 -1711 1304
rect -1745 -1304 -1711 -1288
rect -1625 1288 -1591 1304
rect -1625 -1304 -1591 -1288
rect -1467 1288 -1433 1304
rect -1467 -1304 -1433 -1288
rect -1347 1288 -1313 1304
rect -1347 -1304 -1313 -1288
rect -1189 1288 -1155 1304
rect -1189 -1304 -1155 -1288
rect -1069 1288 -1035 1304
rect -1069 -1304 -1035 -1288
rect -911 1288 -877 1304
rect -911 -1304 -877 -1288
rect -791 1288 -757 1304
rect -791 -1304 -757 -1288
rect -633 1288 -599 1304
rect -633 -1304 -599 -1288
rect -513 1288 -479 1304
rect -513 -1304 -479 -1288
rect -355 1288 -321 1304
rect -355 -1304 -321 -1288
rect -235 1288 -201 1304
rect -235 -1304 -201 -1288
rect -77 1288 -43 1304
rect -77 -1304 -43 -1288
rect 43 1288 77 1304
rect 43 -1304 77 -1288
rect 201 1288 235 1304
rect 201 -1304 235 -1288
rect 321 1288 355 1304
rect 321 -1304 355 -1288
rect 479 1288 513 1304
rect 479 -1304 513 -1288
rect 599 1288 633 1304
rect 599 -1304 633 -1288
rect 757 1288 791 1304
rect 757 -1304 791 -1288
rect 877 1288 911 1304
rect 877 -1304 911 -1288
rect 1035 1288 1069 1304
rect 1035 -1304 1069 -1288
rect 1155 1288 1189 1304
rect 1155 -1304 1189 -1288
rect 1313 1288 1347 1304
rect 1313 -1304 1347 -1288
rect 1433 1288 1467 1304
rect 1433 -1304 1467 -1288
rect 1591 1288 1625 1304
rect 1591 -1304 1625 -1288
rect 1711 1288 1745 1304
rect 1711 -1304 1745 -1288
rect 1869 1288 1903 1304
rect 1869 -1304 1903 -1288
rect 1989 1288 2023 1304
rect 1989 -1304 2023 -1288
rect 2147 1288 2181 1304
rect 2147 -1304 2181 -1288
rect 2267 1288 2301 1304
rect 2267 -1304 2301 -1288
rect 2425 1288 2459 1304
rect 2425 -1304 2459 -1288
rect 2545 1288 2579 1304
rect 2545 -1304 2579 -1288
rect 2703 1288 2737 1304
rect 2703 -1304 2737 -1288
rect -2691 -1381 -2675 -1347
rect -2607 -1381 -2591 -1347
rect -2413 -1381 -2397 -1347
rect -2329 -1381 -2313 -1347
rect -2135 -1381 -2119 -1347
rect -2051 -1381 -2035 -1347
rect -1857 -1381 -1841 -1347
rect -1773 -1381 -1757 -1347
rect -1579 -1381 -1563 -1347
rect -1495 -1381 -1479 -1347
rect -1301 -1381 -1285 -1347
rect -1217 -1381 -1201 -1347
rect -1023 -1381 -1007 -1347
rect -939 -1381 -923 -1347
rect -745 -1381 -729 -1347
rect -661 -1381 -645 -1347
rect -467 -1381 -451 -1347
rect -383 -1381 -367 -1347
rect -189 -1381 -173 -1347
rect -105 -1381 -89 -1347
rect 89 -1381 105 -1347
rect 173 -1381 189 -1347
rect 367 -1381 383 -1347
rect 451 -1381 467 -1347
rect 645 -1381 661 -1347
rect 729 -1381 745 -1347
rect 923 -1381 939 -1347
rect 1007 -1381 1023 -1347
rect 1201 -1381 1217 -1347
rect 1285 -1381 1301 -1347
rect 1479 -1381 1495 -1347
rect 1563 -1381 1579 -1347
rect 1757 -1381 1773 -1347
rect 1841 -1381 1857 -1347
rect 2035 -1381 2051 -1347
rect 2119 -1381 2135 -1347
rect 2313 -1381 2329 -1347
rect 2397 -1381 2413 -1347
rect 2591 -1381 2607 -1347
rect 2675 -1381 2691 -1347
rect -2871 -1485 -2837 -1423
rect 2837 -1485 2871 -1423
rect -2871 -1519 -2775 -1485
rect 2775 -1519 2871 -1485
<< viali >>
rect -2675 1347 -2607 1381
rect -2397 1347 -2329 1381
rect -2119 1347 -2051 1381
rect -1841 1347 -1773 1381
rect -1563 1347 -1495 1381
rect -1285 1347 -1217 1381
rect -1007 1347 -939 1381
rect -729 1347 -661 1381
rect -451 1347 -383 1381
rect -173 1347 -105 1381
rect 105 1347 173 1381
rect 383 1347 451 1381
rect 661 1347 729 1381
rect 939 1347 1007 1381
rect 1217 1347 1285 1381
rect 1495 1347 1563 1381
rect 1773 1347 1841 1381
rect 2051 1347 2119 1381
rect 2329 1347 2397 1381
rect 2607 1347 2675 1381
rect -2737 -1288 -2703 1288
rect -2579 -1288 -2545 1288
rect -2459 -1288 -2425 1288
rect -2301 -1288 -2267 1288
rect -2181 -1288 -2147 1288
rect -2023 -1288 -1989 1288
rect -1903 -1288 -1869 1288
rect -1745 -1288 -1711 1288
rect -1625 -1288 -1591 1288
rect -1467 -1288 -1433 1288
rect -1347 -1288 -1313 1288
rect -1189 -1288 -1155 1288
rect -1069 -1288 -1035 1288
rect -911 -1288 -877 1288
rect -791 -1288 -757 1288
rect -633 -1288 -599 1288
rect -513 -1288 -479 1288
rect -355 -1288 -321 1288
rect -235 -1288 -201 1288
rect -77 -1288 -43 1288
rect 43 -1288 77 1288
rect 201 -1288 235 1288
rect 321 -1288 355 1288
rect 479 -1288 513 1288
rect 599 -1288 633 1288
rect 757 -1288 791 1288
rect 877 -1288 911 1288
rect 1035 -1288 1069 1288
rect 1155 -1288 1189 1288
rect 1313 -1288 1347 1288
rect 1433 -1288 1467 1288
rect 1591 -1288 1625 1288
rect 1711 -1288 1745 1288
rect 1869 -1288 1903 1288
rect 1989 -1288 2023 1288
rect 2147 -1288 2181 1288
rect 2267 -1288 2301 1288
rect 2425 -1288 2459 1288
rect 2545 -1288 2579 1288
rect 2703 -1288 2737 1288
rect -2675 -1381 -2607 -1347
rect -2397 -1381 -2329 -1347
rect -2119 -1381 -2051 -1347
rect -1841 -1381 -1773 -1347
rect -1563 -1381 -1495 -1347
rect -1285 -1381 -1217 -1347
rect -1007 -1381 -939 -1347
rect -729 -1381 -661 -1347
rect -451 -1381 -383 -1347
rect -173 -1381 -105 -1347
rect 105 -1381 173 -1347
rect 383 -1381 451 -1347
rect 661 -1381 729 -1347
rect 939 -1381 1007 -1347
rect 1217 -1381 1285 -1347
rect 1495 -1381 1563 -1347
rect 1773 -1381 1841 -1347
rect 2051 -1381 2119 -1347
rect 2329 -1381 2397 -1347
rect 2607 -1381 2675 -1347
<< metal1 >>
rect -2687 1381 -2595 1387
rect -2687 1347 -2675 1381
rect -2607 1347 -2595 1381
rect -2687 1341 -2595 1347
rect -2409 1381 -2317 1387
rect -2409 1347 -2397 1381
rect -2329 1347 -2317 1381
rect -2409 1341 -2317 1347
rect -2131 1381 -2039 1387
rect -2131 1347 -2119 1381
rect -2051 1347 -2039 1381
rect -2131 1341 -2039 1347
rect -1853 1381 -1761 1387
rect -1853 1347 -1841 1381
rect -1773 1347 -1761 1381
rect -1853 1341 -1761 1347
rect -1575 1381 -1483 1387
rect -1575 1347 -1563 1381
rect -1495 1347 -1483 1381
rect -1575 1341 -1483 1347
rect -1297 1381 -1205 1387
rect -1297 1347 -1285 1381
rect -1217 1347 -1205 1381
rect -1297 1341 -1205 1347
rect -1019 1381 -927 1387
rect -1019 1347 -1007 1381
rect -939 1347 -927 1381
rect -1019 1341 -927 1347
rect -741 1381 -649 1387
rect -741 1347 -729 1381
rect -661 1347 -649 1381
rect -741 1341 -649 1347
rect -463 1381 -371 1387
rect -463 1347 -451 1381
rect -383 1347 -371 1381
rect -463 1341 -371 1347
rect -185 1381 -93 1387
rect -185 1347 -173 1381
rect -105 1347 -93 1381
rect -185 1341 -93 1347
rect 93 1381 185 1387
rect 93 1347 105 1381
rect 173 1347 185 1381
rect 93 1341 185 1347
rect 371 1381 463 1387
rect 371 1347 383 1381
rect 451 1347 463 1381
rect 371 1341 463 1347
rect 649 1381 741 1387
rect 649 1347 661 1381
rect 729 1347 741 1381
rect 649 1341 741 1347
rect 927 1381 1019 1387
rect 927 1347 939 1381
rect 1007 1347 1019 1381
rect 927 1341 1019 1347
rect 1205 1381 1297 1387
rect 1205 1347 1217 1381
rect 1285 1347 1297 1381
rect 1205 1341 1297 1347
rect 1483 1381 1575 1387
rect 1483 1347 1495 1381
rect 1563 1347 1575 1381
rect 1483 1341 1575 1347
rect 1761 1381 1853 1387
rect 1761 1347 1773 1381
rect 1841 1347 1853 1381
rect 1761 1341 1853 1347
rect 2039 1381 2131 1387
rect 2039 1347 2051 1381
rect 2119 1347 2131 1381
rect 2039 1341 2131 1347
rect 2317 1381 2409 1387
rect 2317 1347 2329 1381
rect 2397 1347 2409 1381
rect 2317 1341 2409 1347
rect 2595 1381 2687 1387
rect 2595 1347 2607 1381
rect 2675 1347 2687 1381
rect 2595 1341 2687 1347
rect -2743 1288 -2697 1300
rect -2743 -1288 -2737 1288
rect -2703 -1288 -2697 1288
rect -2743 -1300 -2697 -1288
rect -2585 1288 -2539 1300
rect -2585 -1288 -2579 1288
rect -2545 -1288 -2539 1288
rect -2585 -1300 -2539 -1288
rect -2465 1288 -2419 1300
rect -2465 -1288 -2459 1288
rect -2425 -1288 -2419 1288
rect -2465 -1300 -2419 -1288
rect -2307 1288 -2261 1300
rect -2307 -1288 -2301 1288
rect -2267 -1288 -2261 1288
rect -2307 -1300 -2261 -1288
rect -2187 1288 -2141 1300
rect -2187 -1288 -2181 1288
rect -2147 -1288 -2141 1288
rect -2187 -1300 -2141 -1288
rect -2029 1288 -1983 1300
rect -2029 -1288 -2023 1288
rect -1989 -1288 -1983 1288
rect -2029 -1300 -1983 -1288
rect -1909 1288 -1863 1300
rect -1909 -1288 -1903 1288
rect -1869 -1288 -1863 1288
rect -1909 -1300 -1863 -1288
rect -1751 1288 -1705 1300
rect -1751 -1288 -1745 1288
rect -1711 -1288 -1705 1288
rect -1751 -1300 -1705 -1288
rect -1631 1288 -1585 1300
rect -1631 -1288 -1625 1288
rect -1591 -1288 -1585 1288
rect -1631 -1300 -1585 -1288
rect -1473 1288 -1427 1300
rect -1473 -1288 -1467 1288
rect -1433 -1288 -1427 1288
rect -1473 -1300 -1427 -1288
rect -1353 1288 -1307 1300
rect -1353 -1288 -1347 1288
rect -1313 -1288 -1307 1288
rect -1353 -1300 -1307 -1288
rect -1195 1288 -1149 1300
rect -1195 -1288 -1189 1288
rect -1155 -1288 -1149 1288
rect -1195 -1300 -1149 -1288
rect -1075 1288 -1029 1300
rect -1075 -1288 -1069 1288
rect -1035 -1288 -1029 1288
rect -1075 -1300 -1029 -1288
rect -917 1288 -871 1300
rect -917 -1288 -911 1288
rect -877 -1288 -871 1288
rect -917 -1300 -871 -1288
rect -797 1288 -751 1300
rect -797 -1288 -791 1288
rect -757 -1288 -751 1288
rect -797 -1300 -751 -1288
rect -639 1288 -593 1300
rect -639 -1288 -633 1288
rect -599 -1288 -593 1288
rect -639 -1300 -593 -1288
rect -519 1288 -473 1300
rect -519 -1288 -513 1288
rect -479 -1288 -473 1288
rect -519 -1300 -473 -1288
rect -361 1288 -315 1300
rect -361 -1288 -355 1288
rect -321 -1288 -315 1288
rect -361 -1300 -315 -1288
rect -241 1288 -195 1300
rect -241 -1288 -235 1288
rect -201 -1288 -195 1288
rect -241 -1300 -195 -1288
rect -83 1288 -37 1300
rect -83 -1288 -77 1288
rect -43 -1288 -37 1288
rect -83 -1300 -37 -1288
rect 37 1288 83 1300
rect 37 -1288 43 1288
rect 77 -1288 83 1288
rect 37 -1300 83 -1288
rect 195 1288 241 1300
rect 195 -1288 201 1288
rect 235 -1288 241 1288
rect 195 -1300 241 -1288
rect 315 1288 361 1300
rect 315 -1288 321 1288
rect 355 -1288 361 1288
rect 315 -1300 361 -1288
rect 473 1288 519 1300
rect 473 -1288 479 1288
rect 513 -1288 519 1288
rect 473 -1300 519 -1288
rect 593 1288 639 1300
rect 593 -1288 599 1288
rect 633 -1288 639 1288
rect 593 -1300 639 -1288
rect 751 1288 797 1300
rect 751 -1288 757 1288
rect 791 -1288 797 1288
rect 751 -1300 797 -1288
rect 871 1288 917 1300
rect 871 -1288 877 1288
rect 911 -1288 917 1288
rect 871 -1300 917 -1288
rect 1029 1288 1075 1300
rect 1029 -1288 1035 1288
rect 1069 -1288 1075 1288
rect 1029 -1300 1075 -1288
rect 1149 1288 1195 1300
rect 1149 -1288 1155 1288
rect 1189 -1288 1195 1288
rect 1149 -1300 1195 -1288
rect 1307 1288 1353 1300
rect 1307 -1288 1313 1288
rect 1347 -1288 1353 1288
rect 1307 -1300 1353 -1288
rect 1427 1288 1473 1300
rect 1427 -1288 1433 1288
rect 1467 -1288 1473 1288
rect 1427 -1300 1473 -1288
rect 1585 1288 1631 1300
rect 1585 -1288 1591 1288
rect 1625 -1288 1631 1288
rect 1585 -1300 1631 -1288
rect 1705 1288 1751 1300
rect 1705 -1288 1711 1288
rect 1745 -1288 1751 1288
rect 1705 -1300 1751 -1288
rect 1863 1288 1909 1300
rect 1863 -1288 1869 1288
rect 1903 -1288 1909 1288
rect 1863 -1300 1909 -1288
rect 1983 1288 2029 1300
rect 1983 -1288 1989 1288
rect 2023 -1288 2029 1288
rect 1983 -1300 2029 -1288
rect 2141 1288 2187 1300
rect 2141 -1288 2147 1288
rect 2181 -1288 2187 1288
rect 2141 -1300 2187 -1288
rect 2261 1288 2307 1300
rect 2261 -1288 2267 1288
rect 2301 -1288 2307 1288
rect 2261 -1300 2307 -1288
rect 2419 1288 2465 1300
rect 2419 -1288 2425 1288
rect 2459 -1288 2465 1288
rect 2419 -1300 2465 -1288
rect 2539 1288 2585 1300
rect 2539 -1288 2545 1288
rect 2579 -1288 2585 1288
rect 2539 -1300 2585 -1288
rect 2697 1288 2743 1300
rect 2697 -1288 2703 1288
rect 2737 -1288 2743 1288
rect 2697 -1300 2743 -1288
rect -2687 -1347 -2595 -1341
rect -2687 -1381 -2675 -1347
rect -2607 -1381 -2595 -1347
rect -2687 -1387 -2595 -1381
rect -2409 -1347 -2317 -1341
rect -2409 -1381 -2397 -1347
rect -2329 -1381 -2317 -1347
rect -2409 -1387 -2317 -1381
rect -2131 -1347 -2039 -1341
rect -2131 -1381 -2119 -1347
rect -2051 -1381 -2039 -1347
rect -2131 -1387 -2039 -1381
rect -1853 -1347 -1761 -1341
rect -1853 -1381 -1841 -1347
rect -1773 -1381 -1761 -1347
rect -1853 -1387 -1761 -1381
rect -1575 -1347 -1483 -1341
rect -1575 -1381 -1563 -1347
rect -1495 -1381 -1483 -1347
rect -1575 -1387 -1483 -1381
rect -1297 -1347 -1205 -1341
rect -1297 -1381 -1285 -1347
rect -1217 -1381 -1205 -1347
rect -1297 -1387 -1205 -1381
rect -1019 -1347 -927 -1341
rect -1019 -1381 -1007 -1347
rect -939 -1381 -927 -1347
rect -1019 -1387 -927 -1381
rect -741 -1347 -649 -1341
rect -741 -1381 -729 -1347
rect -661 -1381 -649 -1347
rect -741 -1387 -649 -1381
rect -463 -1347 -371 -1341
rect -463 -1381 -451 -1347
rect -383 -1381 -371 -1347
rect -463 -1387 -371 -1381
rect -185 -1347 -93 -1341
rect -185 -1381 -173 -1347
rect -105 -1381 -93 -1347
rect -185 -1387 -93 -1381
rect 93 -1347 185 -1341
rect 93 -1381 105 -1347
rect 173 -1381 185 -1347
rect 93 -1387 185 -1381
rect 371 -1347 463 -1341
rect 371 -1381 383 -1347
rect 451 -1381 463 -1347
rect 371 -1387 463 -1381
rect 649 -1347 741 -1341
rect 649 -1381 661 -1347
rect 729 -1381 741 -1347
rect 649 -1387 741 -1381
rect 927 -1347 1019 -1341
rect 927 -1381 939 -1347
rect 1007 -1381 1019 -1347
rect 927 -1387 1019 -1381
rect 1205 -1347 1297 -1341
rect 1205 -1381 1217 -1347
rect 1285 -1381 1297 -1347
rect 1205 -1387 1297 -1381
rect 1483 -1347 1575 -1341
rect 1483 -1381 1495 -1347
rect 1563 -1381 1575 -1347
rect 1483 -1387 1575 -1381
rect 1761 -1347 1853 -1341
rect 1761 -1381 1773 -1347
rect 1841 -1381 1853 -1347
rect 1761 -1387 1853 -1381
rect 2039 -1347 2131 -1341
rect 2039 -1381 2051 -1347
rect 2119 -1381 2131 -1347
rect 2039 -1387 2131 -1381
rect 2317 -1347 2409 -1341
rect 2317 -1381 2329 -1347
rect 2397 -1381 2409 -1347
rect 2317 -1387 2409 -1381
rect 2595 -1347 2687 -1341
rect 2595 -1381 2607 -1347
rect 2675 -1381 2687 -1347
rect 2595 -1387 2687 -1381
<< properties >>
string FIXED_BBOX -2854 -1502 2854 1502
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 13 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
