magic
tech sky130A
magscale 1 2
timestamp 1697704145
<< nwell >>
rect -358 -397 358 397
<< mvpmos >>
rect -100 -100 100 100
<< mvpdiff >>
rect -158 88 -100 100
rect -158 -88 -146 88
rect -112 -88 -100 88
rect -158 -100 -100 -88
rect 100 88 158 100
rect 100 -88 112 88
rect 146 -88 158 88
rect 100 -100 158 -88
<< mvpdiffc >>
rect -146 -88 -112 88
rect 112 -88 146 88
<< mvnsubdiff >>
rect -292 319 292 331
rect -292 285 -184 319
rect 184 285 292 319
rect -292 273 292 285
rect -292 223 -234 273
rect -292 -223 -280 223
rect -246 -223 -234 223
rect 234 223 292 273
rect -292 -273 -234 -223
rect 234 -223 246 223
rect 280 -223 292 223
rect 234 -273 292 -223
rect -292 -285 292 -273
rect -292 -319 -184 -285
rect 184 -319 292 -285
rect -292 -331 292 -319
<< mvnsubdiffcont >>
rect -184 285 184 319
rect -280 -223 -246 223
rect 246 -223 280 223
rect -184 -319 184 -285
<< poly >>
rect -100 181 100 197
rect -100 147 -84 181
rect 84 147 100 181
rect -100 100 100 147
rect -100 -147 100 -100
rect -100 -181 -84 -147
rect 84 -181 100 -147
rect -100 -197 100 -181
<< polycont >>
rect -84 147 84 181
rect -84 -181 84 -147
<< locali >>
rect -280 285 -184 319
rect 184 285 280 319
rect -280 223 -246 285
rect 246 223 280 285
rect -100 147 -84 181
rect 84 147 100 181
rect -146 88 -112 104
rect -146 -104 -112 -88
rect 112 88 146 104
rect 112 -104 146 -88
rect -100 -181 -84 -147
rect 84 -181 100 -147
rect -280 -285 -246 -223
rect 246 -285 280 -223
rect -280 -319 -184 -285
rect 184 -319 280 -285
<< viali >>
rect -84 147 84 181
rect -146 -88 -112 88
rect 112 -88 146 88
rect -84 -181 84 -147
<< metal1 >>
rect -96 181 96 187
rect -96 147 -84 181
rect 84 147 96 181
rect -96 141 96 147
rect -152 88 -106 100
rect -152 -88 -146 88
rect -112 -88 -106 88
rect -152 -100 -106 -88
rect 106 88 152 100
rect 106 -88 112 88
rect 146 -88 152 88
rect 106 -100 152 -88
rect -96 -147 96 -141
rect -96 -181 -84 -147
rect 84 -181 96 -147
rect -96 -187 96 -181
<< properties >>
string FIXED_BBOX -263 -302 263 302
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
